`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
J3ZjR78g9U6TW/k7DRm3VqfDzpZ354rwqnsQRw/TZ5l41k1Bg9NTJ0HsS9G9lwfOJcP3luoAq+jD
5rc2igEj6A==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AzT9syKKSZw5rAz9a5JDK+9XhqYc2ZMt2tCBz2q49GoOoxD0a5CUV6je2Ql+S8RE2NZnyNZx6XtG
wyHghKKy4D3x8yzX0OBctKw7s0im3+SimFDtZ+49NXoZ+VIxbjFukiAEvflenrL6d6hIfxq1P3IP
FRVPrXrCevbNYCQeEvw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZLV8A8YWQ15MxV3M1skf9KnbFuRaNq4IZvXBFFNi4HXjv4PZBn2w+bzKJSFXybOoHcZ9s/3ovI98
n5ory8+rjBkp6YFvOiLN1z26u6tNjuWSBQU8Bqg/Z31KBpxyGxRlZLaMJEwC3PDhAW8MeWLZhvqy
qsVBQo+evb9GVmtKCQzsinqjBZwDMgrZQzW40NSF6w7tmLGXqm/kKzbYIFTnT9JlCoxs5eESxAEp
dOA4MdcUyGUE/MSDyDaPGu7KAd7Ef98fRZQ3MFyyaiTpCplspF0GK+t/R26Htybe2nYCb2QdAn86
pj5HZrChlfaLJiXR60XvdB7CGCH9+Te79rBkqw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oxG9OxvuLL507gQTO27sMBhkCbaIcbL81Lqnx5DFGwrx75ZE1DabaxKIscU4UeZljrmXX1MgQJ3c
sUv1je6aAN/DF/OLhpZU/GcjSTzmLaPxE0r2Q+d6hh/0fpfeUknGehb44O+AsIPSc8eglo9hZJps
98DOdlk24o+IUsZp/37VM8WV6LUOoqZ0kiJmqc68B+11N6ql4QvHLYbkFIh5M9FeX6xAlw/GHZJz
TFnTsHSIlF4sQ37bo+ozTAUkmu9SO4khaHTVB/eCZp6rxp8/wCwknte5qQMpeGlfxFiZdoOo6ysE
VVHZmMfMrLVknyN8ZgBL1ksSpfB1dp731ghn6A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sQaTKq8sb9ucuzMqe0gZMJZuNsMqFGq/fYgAyFoC5kE+n1HGlTxX7KEpTBsggn3qCUVFh+j2MgBj
84eQ+UFV6iU/vHvwSZY1oK5v4C9GQiDbZHM0LdXhTBioSJthIg0oRUb9QwHz1Yn0dhV/alWV0eM7
sLSTTKWjmfdo11/kLflR7vtwAD13T0Pn6GX6PEFI7i6239o6o8ZpxljESkuu9ThpX2SFHrFfifLy
IF/zqB62h9f34jCu2f0EpM8V/4ZgMjO+wT7jzd9L1yhyCLkN/U3gA3usDP16xEDpfEXw9Hm8HD3F
bIB/Yeg4MOHZVPjaWWZ64fdoxDzBkvfMWTTZ1Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NDaDpnP23TbnRd8GBgBvdkK7cBv7n2lhI/dKbVeUM7bx+c7ewW5di+guGvVBmT258ypt/UzQSK/c
vkdCMTs5C52dWr7mRa330cw05WJlyJzbIgRkGxz94l5gmk/5EdNr2FBX+mEVYxbZUOtdRgZECsL8
xZcrVb8B/anXbPkfPKc=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mZD80mh9jOJwoWc0TyMSnXzNGQKlg5nEp++zY0RfQ6JkDEGAq9bKa8VcsKpnVdJAOVUl6vec3c7s
NPa3FIMBNCq+IrAhNkD83TgdEmFyfxUgi7Dc0pUqH8LeVXsg4GRQqRuzDFn7N9YTALnfA0Z/pDn0
Aho64FtbEyyn+D0jYXuMhsFD6RjUsgH67tX35eAbMDxFlEKM/9pyMxiNqTaZw0HGnAPEEtfODJSx
yzw64lC6/xm1gZvJAGhIoZ/dYaQ8uXIfnpce9ei3YhflOLM3f1U822doqSrjAvc3A6inPE2dv9da
0PIRjnhIzS2V5olqAc0Me93P1n6O+DV/3/+AQw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175280)
`protect data_block
5vQjzbIKvdRYPs8u/Z9AV8lG2x1T4+qT3G6Ui4FvuI7kdTzI9MUtKeB2W88nbXAhHnr8J34CyuSj
nLfAket8gEXbXpx4XL38axUfhfrUVlxbLBznNmIol3Qln3PwPx7zeArqjpTwC/CCjb3GDMxUZLlO
mFRTPc8gXUhe7yerya2h1yEGazmsVIRvIDb19ISkjUzwIfzTdPxkY8gyps9yfiWBemB+PU4mj60Y
ECQa5Bb/Pp1qTrkiTqMUr33AgP+Ip0ER9TAU0/imWYq9C94Fotbwr6aUwmnKB6M/UBukOGWt6PEf
/oH7X1XcV9LW9vcQlhtd0kXU4j+oCMBVc8utO1mWggedX8a47UXOQ/nJWDnh4yPER/YHxhjYhp/V
jM16QXJ480MBB5gGcVkv+VL8fwBPqN5p0O560N9no7rf6evtBAwMYLU8UF9l1bGQjjOcJdp9+PJO
GoBEQBLDAZFOPSmGH5sw5/fWDz2XQr+PjV6GKj1ZsD0npopyLISkBxWnyNij3zU6sYJegI4Czt3f
kxvxEaCvkRWFJcMovt8I9rRr9/m1DXVbC4M0A0xhwt0HcQ5J9RDMTRlzXCmSni9FlIfv4Ce6VxcR
QeYrTUzL+qf91hU/ieGaYgnl4FifvAmXb8Zd7xf68AeRMHqIxvl7bUTQ40Rv3QH8eweODX9CelWy
JrD3EkOcTuG4UcMugZVexsb7cDQOMGa4PESe46cwP+SUhGTYram//EKYOkihA9DR1YQ8hlnvvdcQ
+IDBXpqXJm1FVmjaCuVUfrlRtSYE49G/fI9fYnG6zu4YzJ+UfV4Q4CD1X/1D6NGXS7bY9rTroVUK
l6/Seb2+jWcvm27c2J2DgTjdty3mXfMnrYhKpoUIYjxY6wvcvcwylaK9IDnj+ZQVTrTGYF9dIjHx
C1T2NHk76kyjkNDOxwKxo34kYLnyihSAfEiLvNhpry7nREmP/VRFMVHEEnP8TnoIqQM9sMjCrgSw
3JxuTZAshagM3wfPXRq77OFCqNU1T6cBnTRSbDQ5T+Ny1JagX4rlQBCeOtHKJMYmiB0EMOZhmvqo
9liKTaU3U3EMOb0Le5LkVJJ7bVmKrAQ8xjIeBK0mPW2JuKd6i211vCQFLkKUqOmNVeS0pQnpljLO
+++bOVdQ1NmYyRB0SqjofGLtPKqHAMpsIzLluloB1djSUfHTmSkhx33c0pDPb6i7A/8n624KqXW5
o/1DZH8/6QjTJxqRzRgStdaE0QA60dXsaP30SRmJV2Z7nQjmhW16roRB0tsskm22UIKCUXf/fuPE
l3ta8kFHuqgV7ORwMQC8RSARloPpqnWPC8uzKugdAZgDErWKIlEvbDIKqI/hnD/B/I9yHkoebfyd
WrFZWzkoyuFR0PCS8jZQSzdhRuskT0mNAyVAT9z27z0b6dYYHLf7oOveHxIAN2+UQY+EcM5B3qjr
aYOTtDaXCS2wV8uebNJ79MAM1EV3bj4uZKHAMoWRyGTIdTdRmNmgZ+u2gk8FlfsIxxNZ4rn/Ky2O
BGjnyABeQeuG8NBCwfgC8mSResq8oxajJp4UisGpuOvdp05csxao1imAFhjLqevO2KYlgkLHM9Pr
yMnbI68HXVXmvW6F0xz9XWD8L3+PSkcjIhs99xO71DDi8E5pHM5UNpMxssRW1NzUseafIObDxIoQ
Dm+HuyZP1tjYMYgOzr7qGa5IU9Jyws/yA14d/AhtAfihALO9zvyuDh9oiyKS3k0OqiD+g8wojicq
Cx+rwRVRX9xYMoYyAEznRAsxr0v7mo8E3y1rcGH3GReir91ZswjLTjEX87k37LolUxE701fDGsW6
SEinnHDMZOPT04odxuI3TszUYC8aIKsvGONkJ4olHclt0pO5ZWAnevEJLIiM9RvtOpDnAcgm75/e
RFrlBYeEmI/T5pVQ1re02p576Eiv6LJSvGPE7NyLGxIznKWsB0StLTyxMx1CV8E+c6SbnZUdMlGa
67/R/vqe4QhRr6/BlPsDgmVM6rXdHt6OGCscohrzJEZuqA0by0D/nlRRV5Y4itp2noSzJD2UZIu8
piQswZImRws3VF3FtJTY2ZYO/XCHGrkcOb7+7bFvquysYw9f3z+MCriRmxbUrxmZNrQjAm//h+CD
h7yjZkkOSHS+CfaDabW7OPciRz5KWJY9HOwmGyINmoruIC1xrIr9Isb5K7vmspAB2A5aa4qiGlor
tiG6Kq/dpBWqRhy95wcKQo4Hah70GxxcrqsaAoNdypLPcdDU4HC/DeF+rxEtU2Eq+4jD6oGQl4vf
cAWj13HiJk0hoxcjYsTi0QkPyV516/mrehWK7HlnoKQjYMgWKST77XNcdtM70niYXsTnniqxxBrO
6G7L5elxvCKya4z95oBbVoZanwGFGra989lV0kFXo1b+lucTghIrkp9OKhWYubEwx7lg3yhYQwLc
+zUv9kGI+2QcQppszWsDPl7zFDoYTahFrJY0rUBHabyoKgapOIzvZeVnQHqr1O//qY8164F+Jzca
BsbYFLpyCSHki+IwDh9r/7V/L1D11BLTydCEJCwO9hHBQ/KN2rDGDymV8A2Jd4a6m/O5ncpJ0RKR
O7MPTY/WYIL7dvruxa/gJevQZHP90iZkcuOW2t6KUhkMcCIjsu3q9FQiBD1aTHy/vSTiVsnTZ5UI
CdIWkWgIGLJT2Fzx9A1UhjZP9TdtScBr0wWDLTx1Aj3ug0WGwvkt6khFw7WcTZuR2Us9xY/HeKjD
bQQzvPumrUZq/f/L3Lh6gcZoSC7Z0LCiRWLuQBZV2F3/FJd146pPlpQEHS0HzZzQXyl2/kjL6r/F
FsnOyaCcd4U5/9SfLr6La0Hjjfb314iHD4LdCz/hPmtQwslNt1HP7lt98ZqS1dh68cC9aD1VEy1T
r0XKiP56xexJHliIMSLHfwOLFuUHX0c+9CAQ4mzDPVP4qQVimJXyhzlUKz/cnNqB+gdotof8bY2Z
dggYgs5aFy2g5i9a+Aq9vcfzGznabAq8XmhvHp3iP+RVKTxckcAq2bqBSUqM19KmHGGn6eYhcDPA
B6HH67Q1gkxGUMb0kYZlfXSDRC/UeaYWG5SpNcvClfecjL6cJLuvm2bdJO67PEOhCbjK0xaJKyGR
zoSbpIZYEtSqv8eCZp/5XD9QdCxbkYkkXNmz5u0tpQaCZkyrvmF2XjvYmmDvL+hIRsSiwI+q074K
Z2fP3EXqhrFdqfVeMb7/NN9hubMFWdvEOS2gjnNKIitzgKrIkKWPPKA8+n4e+qa4/veRV2n7LxMF
slg/R6KwK4TptJuwz9Z/7ZNJh0Ct9y1rfNBqej3vxxfvtjhTk5emyI/j1iGMTulW1f9XDGiTEb4r
VU32CItsH8pc1Y6nPpzGYuYn3vItQ/aIzlK9Jy8rnoocxhEb6+v712F2J5TcixeyrUJhQ9+7C5+0
Hvb+OJBvImXNhz8rS9sS178ov5YzBH7d2zeElYUuML+U9NMSSvEMgrgfe3GmN/Kf2ICkwuB68lwv
mai/hplR8lGRRIYp9TZZb/Q59/hKKMR687s2xvGxPaFhzA/piu2kRj3LLQdyiomPWv6W/opEfm8Z
VjUK0w0TSv73x1csPYYND2/ujsCYvfPlKjcohrEM+g8mw1ncMfWZNaYhxHngLPGf7fTyedDlGXQt
seFEqIzEQuqiH4rvf2mxlz0Dylls77lD+OZVfeWKOwX5igi/bdPebEWvRPzXbFryXydVTl5SJ3jc
BECOoAd9luztz10kPotTW8PTtBstmOhDcaHckFksCtgfs8qlzR+XiTVjKDChkJMusXYJY9D4XwBp
aUBedspJFlJRCnuY2Mmdc+R37a4PY6Y5iOeLWVeb+3o4C5Xu6Px8gzWqtQsPiQrWjbQvnrg+iDEM
1mfnyWhGMGsxjUEewemCzPgJlcGcCmSLqP5P1VjCnjMcGutrQYGwShyalA8Il5IoaG0azc7VvJjM
6AIkBm1kVXPu6PujyfXmkY2VX1ipIrL28xj9T8q5QgmReSSxVei1/Qot0T0d9vwo60gEP9PoLEY4
BLRsHQAt//b2u4b1SYf9fa9iwhd/2Bdc39Xr3Iq5tNpQXgXDlqilYJytkoNlUnKG36Cf2iFelGpk
yrPX54g127I8McDFmqo56RJBcnfRe7D7qg8SWfaQr9gWWC4pkyTVjM7hjd2ijQSfaLU/V4SbSuAQ
yHOnGsd+PYgWvy3PrqtTPu4GqQVS6PGCb/FKTjlWeE0PYnJUXUdGSIoRp06AjIFQ/WiKWMZwBjs/
rXl0inkihjNyt7Qr7Kt0yxaAcTffgNh2VKRpw+/CKnu6gIhTDsIJhdUHTz++wPu6xvw4ZBR4SAMd
/tQ0gvd+7vRZ547oRb6fNDR6iiHZpMEJ6Bnu3NTNkiug+0Z9dX+aKDXTyqqczcraxQ+FlBaLFGn4
A1IePz97Qnw6mP8LB6Vo403Z9i3meOxZMmWdUuU8hcqdWrXWPwAfQJNngTfmFQuKU3S14pbCFA38
bZbKrVXyvKOygS0BulMHm66yF7DItFdOaEgRHDbyryxDRcJYJ1XVsZ6km7K9usF2TD8z2ZBuPixK
Mv5tQgWj+rl6ozjbrzTbJY5jwGrA8+i16XSLQf1jodGeHfKIVQyL8RURwHrqA+ONoKJlz0TrqlSl
ltRGr7AsAc41/y2bTCv7FWB7ApVlFkHDdE1N8gvyh+2f9In7EpyCo5kpRo3DzsSfhmbAW5gK4Tiz
xNbD1a4FnYVyubJEaLJEgIM5EY6jBXGYZrEYW2n9O4l+M4flbwOMSwNEsUo/VFXIAn1Bu+83c0e8
YT2nAlkkYgNgeeh3E04Md9ci7Bqb6KrR0wYyocHYV1ESA2Ufr7Hzx52BKengVdm4ZkwIwTHHVbcm
5Gdv3uDCezB2LD8zk0ojxvTIFxEanwXPSyzWX1K9as9bU+HK3RT0P8pDmu6ycBWhnvdgmluKQk5P
kG76v7mUeToxQZm5JC9uaOnDSi+OsnVYYQj6Q0NgURYQYZv5dB6qSUSM42h0Y8hwx1YAK0tWt21y
OVpS8THXWWGJbwDvW+vZ33LoASQI6EwiKzsTg2RaNqoKVwdPIoZ/u9gEN8xWTyz09J77m/Ak3YhO
faJzkWTUzEtLHhelWuzLuONxXjOhA6h2NpAMDTuR/Hb69U6Z3KzuZB883RMdyhO7wLdDUuSANMRe
xZQIcBk3d8ivi/bOz0820geGOHCtPvBM8Oun868qcXgxKiKDA7avf4b5q/esVx2D6XhacPNxgdDE
ivZBbiIdM3jx0s7/8UTLnAyxe+SUoVDkHdbESB22uJ6Sc3S4WggKHrLCvVpuHurkEsnh0c5gftnF
kxOOj5Mmesnfb9ySnTrU8Bmj/TO3kEZAwBZPNrYStPGHwaWCFqjE3TVOd01rlbNxJe2JIQY9fIKD
ALQjqvh7JDkdtKWT2nnF/9s3Kj5gWqX6uvHGKApbnpmDGQGSSOoXz7LMdM43umksLQsja/lFgrk2
rH2LCJ/AZo9tEWJ3TRBZ/F9hYda8QsZqygLQbxn9C83qelQG+ShT+qNxMu4ZcCqnsmJkDzQJZs8p
NfXmitrihjMtUKR5Qmd2I4fomJ5nkCg9VOZGOmyE9yiT9sL6/oqcfLZnhEG5WHUJ3xJu6jrCavLY
Z+ZXM/k5AYn07LTMQ2DkbV+hOc3kmxWs6Uh0kmskZu3xhqkSmVZmRQuChAahzj7i6oU+g647iGfp
fiHos7eYGxEpKdRr5XsfFPyRImzWzrsylg12AFQ+agPJMqLDYT8iRpIfTRK6SfX64HlODNUkHLo1
f0nxrPnIOA5pO/hGeDQ15X8kpR9Ci60gZ3ji4/sK6Bs2HVfLV83YGFUE2bnGKmTIDmvVwg+yd4Zv
tBU1RonMrw9ZOIrTDJikeeygJPtxb4MeY74rGsZkkqH7/f0VFF6fEMtgULjpyKBeZOg46WVOtlj1
vHG+S2ium336Cdi6tvoqC1KUOEZL389OMVQPZbGK5uoqnRXO2J4k3K9/32UjzUNxiuAH8PTYrEcC
YnkQiOGv9p9rveFhTBJNiZK4x8/BKhBh8SRVPtKGMlM5D+jUvEYMgh+NGJ1dYPdj4fm0pp3KrYG7
dhWge0P1EZ1o/W4Alak5cSx/l22aQqfXaSPLwCbmaAx8ZrgmqIJajV2fassT0CbYhkZabEnn76Yj
d4w7vHe3GHqu0l15mBJnlvayjIN8MrgxE+5CRcb0nw7XmYkivpv13efmsX6PXE2KPw8MYGxgVaYm
iYWMMH6fwHzILi6nOU0p7HjKH9pD16SPX0CX2Iuk4ixyyUJVMpBWlv6V9XIhTHewjyE+YTPE/Cz2
2qXyLOGDTPYmUhoBPymo4AB1cVG01SdquuZ5kCL7GcM80jkDFJnvfEX/IM252fPhNOOTl4u5vidd
xPp65K0EuiUTcp1UP/IgJabeMor5O2XkC9PzuAbl8GL05PDZzkqehO2nEAJ2+yInqJa3zwIgat7L
9o/B9ToyNWAKjfiADO+sNwbEuse4P9O/R9P3BL8GUzSO1rQZqJwZZXPjFxPIlETl9XOaONv0q64S
Rrn0VBLb5NG2v8FlnCbPmool7rR4N+YhqAknSkZ9SN8fdinyf0yMDvUyQ57HL+Nz7doIrueSGi5v
kGYos8Zc0wgj0snElbqriAE5khGiFUKmU7C9Nb8ozmd09IZ5F4663XcGR4UAVfwGts+QigMLnpfk
t05HedAM4T3px76EspqP8yNbQ1tc/EQJ9/lfmqTkoQyBrcdt+TKlJmdmG1uo7/stNef68Yo7emrl
wOB0hES90jycpJra2PlUZgluaANofjnhZnh0OmB7vUW/9CUb57B2S/b4quuA82eMS+DrfTG1gRj0
tyx7WLd2LjDdqIKo9WBhEcUV0MqfcSALdJavTmKXKbFRcSmWFCL8RepnyIAOxY/8FoUN6ww4KiMF
ppFP/mGUcDScreCT4rs6tsbTmYV5RKPhOGsirQpaQshH1gdSt3fZAB7qmSBD8xUHDks/ArnLyn7p
xkkfKfPmUxYE3z4mC1mstaA7olKPriEjILTBbYP7Wg67+dXGe+/C6C3fz7I2B9ogssCyepVj4ONI
ntHts5I6TJoFF0mLMF7wa/X4ahg1YflAXgfEAVLfBq1kVK2iAM+Pj3l2fnBbFxUcB4PrYQGY8o3e
2l/SL8IVG15CBc+9kttdZzlXV4RHw2BB9GKBsQmkGqSrXmoxnjRhFOOe7HMF74WqSoKw3Yh8mioc
zR4M57m9+GdYRY/P8+fVrJoChspSEq3RIubdN6AJ2R5NT1+VWPPzmJJbig2MKdJAlCe77lsOlm2U
rQI/ppLYcJGfgXkiVldlh6WWsdEl/aVQjJeqRUT1+bGGzxPG+wuj9xQ/0Gs1dMqFreqZ3Fc0Pr9g
RTL9bCcuXwoKilU3pfoCkKHMAkOjFEZmlDKqUG5BLm9Jon9Xh5ULcmKuPnPCP79q4EWhZqjpjzoL
FFy2FhSHZz/ZFKl9v6X3PF0hTSrAafc0fcqUhaAyIK2j0JbGvcgmVu/n5OabyfGDPwwh2XBzxPSn
qSJ0KkoP0rlnii+Vv7LIUiwmM7qS8QddtMQxlaMIEW+qHwLLAFL6wSihmOvxb+iH5rJvF4TkPQ/D
RpAP02Y+IJk8hbTzOQlaqd4wG/SkUcbQ6AhSApX3UuVpr6QbVdMK2mSKwFDJeKf9TZYGgLkAtUhH
ygFWV0gGHMAMeXmPgBMUlBEsvOY54m2GQ/yH8iaQEnDaNfsP5zAcRM/IswQ9EjuFbR+07Bk2M5TF
4C9MJk3Qk1mct8jHDONmVzSib9ENsxUJKLJuwyFrELBqI5MG0WcMunHN2DiAhR2FkxqbzrLq0Qdk
a9LxzJtjPCUDKjKaeZk6ALN8p1J51Sz0pC0Ey+geXsXnH87ta2qtcG2VpCW9G1ZJjkqNv2TtcVw6
+8ZW4IUmCzLY7HRevQ3RP1l9kW/esdKx/NTY2yQzKmToBQ9BUDJsn0YLjTbSP2uWTFGGL9v7eQMC
AFPFx31fp5yUng/HQBaNS559NSsaOHTsDGpDlpIFHOGX5+6cK9atc4L9kvkD4np6nFEhVW1A/NOW
bvcOOONp2qmWtiXqmt0GbKxS6DKXjm6Gad8lz0niQZc4jVCJTzIoybVJm6VZLs2EM4ShZsgE9kjD
5SpnU4I2Ci/TbkgrRrbbJOoDywX40F699U9Af0kYyXx5MMwG2jywMFNG6pVcCkMucATqHio6yKzA
tnkZB21oGZCZ2dff/amrFBY7k15x7PBHQZE6Bum04CKcE7I8ZBQWtQh2OUJVJcrSdHLIubKv3lU6
YBlWDixLAXk2658KHDEBI3PlPDKKmaTZYDlmqCrkCnxXoD7ZnPYnyUoeSAuWUlDt1DrmQmnUPLyO
aPlgJcXJb06rcsWVjBne8Lld8ZJPQLSY+Jn+OgNRDw/w4GRFL9JbEypKUIasK5rQsYfzw8J+T8Tv
G+Q0pbNCO/rjzcXqW7ytz8teP/pz69eDQyU6l+g/Skwuvh79m4SUgc4khXNUOiqBNOKNmgW33ZkM
+xBx+riw68phwTZzXm/UemDRHpDULUS0BB+srtQ5zdXWKHKWEVZvZEnUPUaYPg+Cv+9VvuI0Llzw
wPMsinAt0TgjrDXoGIHf3+OC4eaT1gsCGD2dGNun5WidfFnPBjURHq3kjjUT5OiIqEfIQTDNGcLl
AfI/luLuWE/+k4WDjPG5JVWz7xtrOGzQCX0VgTuY0tSgn0d54nAs2Rut+tajDR3bByasnYxaVbmA
oZOLI57f8xLz+fIhzl7FhJKSpC2O/AadqE0PObG8bIFvnDD/EjlHIHumlwok+xrl6lvPob8gAuqu
SBkg3AiE7uL1SwXYisNSvFIeGE6uqGN+WUtDCx3/9k31pMeRr0YYYpDltTljbiAeha5u4/wksEdL
UkPUtjV/dEvILv2hIH3Rrux9UUM1Mfdro6eetHrJZqD1+gokfL2Y+BAgnZjAMHwKR7RQYRwzqp9N
S6r31zTq8tkndXbWdzzBILWU+U7t1kPKwfQgXKM2zbThy30/oHdRg7ZDDAvq6NJH5w4LrolzLjKy
ma5KOKFxTa4VZc9PP6JWxCxwB0WsKmjZ9gypSKZ5W/14vltsAWm1wcsz9ULCN/HuCi8cfBgMeGGm
uWE8Uje1z457tbqeqLAI7SJIJ4C0KIT9KYSf7dGcXfGFU6LLK0QH29vRDw62c4fNSERL1zXYjl5E
7Zokzodtty/9RdWHqjVjqL98OBRMNvotZqToJ5DSbmXfGiTQNeMq0qGJNJmmIxdDzP6U5SV8eWVH
WxsLJ70uu1oxfT//9xUrElW/1zvQfXIB0NVoAOA9sdP6I9akWf2YBB7CeJgypVOxAKOetp16PsSU
G/PA1eZ7GntWhLXT4s7KYkiHXB1xaruNXJ74PDSE1gsCnciZ68CnEbyPANLskdsxOk/MfjbXAmDz
Wtrz+Bi8xeQOYxnMLKLbUdlg4z4UaCFokoASYVGji0r6jb2Rb7jcBaP46wmnPGVkMNAkRSOGxTcs
Iq6e1mT4oO/8K5oF4J7XUd/2pT7nxa6YZk5DB7UVUXYyt7m934LCHrwVuUB+NvIgRDEogm7HYXoA
OsDwwu6WoI9pStKj7Xet8Of+kBANulhMeAbh+KnxklTa9DWQ5115w6iUflpZV8PjhbREFS2Eu9aJ
qQPfh7ft4gHVmK89fY0qJce+sv5h/DhhAqelg7ED3Xb7wg/jtAPzmOck1EwiQ4kIzXy7FeJVCdwX
tBOJ149Yu3oDtTe7szIO2Va28n/c1GIJtGyxakHIC+OeITuMdXnx/Sfl9j8PKnBTihV5zjaybpTV
3MtJC9SCFxcd7UE/gEbUMqw7vv/TPB5gqJ9s7fyuIS2mlDaiCano/teVlBiA5dccn4zXrF1pHAtv
m8ZOX0QV2UbV/6hdBekVybU1oMLRSRj+smEtU5fEIaRpiaFO3RlKZBUmv5SYc6JrrzPs0yRsKDRR
52P2P6lel3geNwpTVybK4e4YIvqaFN8y1aa397hcwjrGZn2U06foJkrv9aMnXFKSm6RzgE8sjN5B
e1GtS2QgF+qviEqvv16sddnuXSmHIEAVEybKFBAAqN1r53wVV7o5Io+Aa671A3GnQ7FFOt+dl2UM
fbrt+On+3cL4hQqMgm2lqQJ0Z09G1EgGuOzZWZn9uuAX5sz1PWYWn+peqv/9ez9DxsrBuobrgphV
9vLOmiAg9YPfXKmVsHrw7BF1zrojdrcEOrSkbyuUk4muOdYs+uZ+OwWO+8YpFIS2HSjziBMyZ1v4
g/wzeJW4cFdSOM44RyEP0+EwtDXpgf24RqlnOpWzpRrbbm+G1/2gRrllcDSbvxzWoeay1G302/A3
1K+Eosvq882FdMCC149kVfTsSaRcE6HWg/0jKtc3l+QTB1e8cJ/hghlOteq5WGmjLLNh7uzNP6U9
mMW85ooCCB6PBj2zg/bcVO1OlGIWUUzN4kskrR5jQE013EFYh6uZ/9ut2bxMIGe5KP86t0sybYCA
k13eh9/E0GPCgBtBcBEqafBkMeKblAaS9AlnUjOAAYCs+zGw5+NrFzLhmrjJ6gehwrYx5vm5vZKB
FKs3TkQp+ED4WVaKEEugDVDe56JoAFGQBRpz4umlIyQC0DSf3rLXJnRhlk/no0ctj2xOufxMOnew
IHiqFOOOTUnCKVqTI13r4AQTMTOykpb1TbXLRaaQFs8gjTxP7t/bPWI2UiXp1V0Fw3Jkd5bqpAEX
icUQK83e90uGQQCfJoJ7iMMFgulTT3dwEdthRqXs5ezp9yQnaKyZ4mmVo06fP9FU+qMtxhFBeP2m
FtRpI9UAyv9wuz4Nfdp+ABy9NII770jIOIMdXvIkPvD19xsvGTsbeXV5K4UhINHLuENkGao0UWtj
RaeqavpFd2EEOVjKe9Hxvl+d8lpMEWdqRkIbwSRhEN5X06/vzg/nQRD+6qkhjWkYELR5r9NZgfJd
0Tou4jYTPQ9yNNjUNDnZo4I0XpVqCjDwc7JK9Rbz1Ww3HxHTXGwMWI+c1nflTHZ7DL3+/zssdH8M
nTVrN/fbWQDiZ6doOuZJN1F5d3KnXOzACxa8FHo4N6ozfoqWDkg4od6ZdJcYZ3ZWxP1V6ZTALvK6
wl9NhdksYmYYwGQEmnPFtx+tEcDTKgI0OwLpNb/nNj2RxVBAfQSE7rAI35W1FKVs8MESBZZIEiwE
IcdiK8ibtokjeKdBSm5UwipKO4oo1Oz1XdeekbmxISlN0emI9xnlJskXzpF2pYrkACpP3ci2qJV8
3puqgXFetYg0V1YPb9bNwOde2TZPH19HhOUD/FBFwzrn55OSzjjmjZTasYfUsw8kupAmTE1En/Oy
EFURK65I6LGiwkrYQfT3JVrpGadmdYQFkOY0YSRoZSkqscJ8HC+mehoZjZ48heeaoKjgaBudLVGm
faQz38q30Bseyar1wvZhBGTzMQkmCf74lE6C0DSBz7/wgctvc+PhYfi6r8eiwrtE2Q3yFPl0MUzu
154Dg6oAUmwqAvWCnTYgkkeDgch8U6dyy9BqyZfovzIEXhxGoZ5jzrg1lhXLKZg4ekEUBa0DBihk
rsgmZG97t5u7YN2yKMrdotrlByosB2cUiEflam9oWBSpA+6GZloYo1ufq5tqhSG7eSf1uOZ4ayGC
+SfwIIHH3GERbl6coB6r9IWn5AUnVCbmr3lZ7HqPf63n0Rwhvwz5I0TYAsoRK11z6mRKf1Kurclz
VcEgFMbk8ePih15cv8iiY4fa8A3+G/t3dpXyKX1vneHLjgF03sZKBVm6z0UaHESUwTLlgqZZSKU1
35urFIMNudgBmjkkUZWCYpT4XNxjSs6WvVzR1BIuuPY7cQn1v71+k0t8BSmEuxwMilo/vRaxzs+U
i4qhNR+GPkHgEI9VXgyZVu0i9kyvHxjXJctvZPQPXVY6YrHMoAdsvJSMY34lzFSzniC11T3eiigC
bsj/ZGOi11iaonAgzYCdJRz7Fn/BQ2Y3RTHfktCPV6Pqq4ilIiEbTjKi8i+x/++TQ96RCBxyAf7E
ST0hjKXGa4O67svdE4/g1tolOGFrlVQDMCPmKHBbGeQK/xKfr1j3x+S6lmbrfdYJ2h5ngIo17hCu
lZUOpQ6o9T2xd6R/RWoW0iVAg/3HJvN6fKcaUBsaf8I9XVWnQjsp2zn3vAjtB2lIQSs4YKNJYkfH
6LsWdjbe2prQx8SqRIqZwcZQt0EmNOv+YNGYr/ceZLEVKYGVFkwCds34UQBGnLZ7HKPTl4kI+ZyR
75l/e6hkeOh9KspZ/3cTn/fkoKVpncaNyWx6tMN6rcR0YNDz7YXml7VSnLTsh1IHNbQmp8YKf/gQ
l+0brM2xjWoRsqWIqjBOrTc/j1oE5FPUvZSdYli3wt3RotJN6eS8ndgn2ghVqTGH5ekxhpSEOL0d
QerJscj7BndkcoISbmPvrtBvkB041979ULKupvhDq5iRQxaWoljbHWHnv/sCe93drshfoDQNQ4IB
VYi7aklzcXcDJClRIyVudlR8Bie/sGHUUr+CrgEBvWTj1HgiMHy+42ELPWGrgY1uRXkyIBRi+1kP
Jv4OnNbb6zG/dAPVbs6fgFuHLyhHqK3EJu28WIRWSxmN2NJP09DiBuom1Bv9xIsufnG6Pzk+QZMP
v+5w70OAyTtvuw+HZDvSnFOlyABUqq+NHsif6RVuHj+Iy5zo2ffHPIGUp/NHdY37/reiy5YqdB/h
OJhnXXJWi+QoYQKj2ZpGb5OyuQklDI4X5MsYiCneKR6z54VIIVq3nmPwhYEZ51Fn8gG6Dqp0XfPI
Xs+pWwN8uwHnw79Trc6aSsEt2LXZR+tlTk0aIxbl6BDmZoUhBdj/ufyr79ud759+7xmuN+a/OQiT
ad/06Ekujp0cq7Id23fQTV2yMol/ZOoQz+ZkrsZWmfFWNsopmQYtnYa/V+azjxHLrJc9vabyzVo2
axgCWPkOJNhA/FjB2WxL1G8X+Zvn/W+B0um3GUUljGqG4AT05KNHKaycxFUx2LQ6u2gmXr2FvTS3
P7m/krI4fDok6e+/0fYasIHCBlqYh2KUqT0tCABjkzD7k4XgYPuXHaV8BTGRNshqbEFugL/VDTOG
VhYSapYtSEcZydAjY0Zs4VHl0LaaNSklBIcvtnT1UmZLgxTsnCiCFAPgYVhq4vpM3IoDB0b+a2ID
pWLg3+XtuvRRNp4VyfEO//d8jq4zxvvmO5uCBMfgxFu2enEoDuJQG13FtRZUImdXvk/M1yc7IS+A
G2hjqxBJgtabCHiKi9+M9zzviXzScBC8jJ6X8ILmtRr5RhTKm5SIBGPSBWeDQKIlVJMZSgt2z786
sdLCZYm7fD4Vou7Ixzoron26D3capRUJ/CC4IeGLlQY+oTIW6spFmdlQcG4So0FFF7HvJzi+l0Rw
MhnItLgiysYQwQVAqsoHGKP1zuFOeKZrb9bCuN2njFZ+ClcSZfB7K8dfn0jhUn+HcpmQygPFQtcX
S5hOk01MMrExmTf8zHgxSQRQ5rUDrZO6lO/JGY7rfwQnO05VmeDnMW7JoZpBI76d0Qv1Chhs3dHd
JJzfjFpQUdMRpavTgslaD0QUyVP1/rQ99AeQ37atmfz/Jvf/pDCMCowizcxQ9eDmPLH/g8ZVIoUR
HTEV6PpgVoABl/uNWFHsll0PaktF0HmtN+U/9ZtZlFeImMluFkQs3oI11Li0cOaEda1HOeEg7Oya
zgoGfoKIBlPdS7odJ6E+Cj46/jZMfrP9qBJGOEqFV1OpHqc+ZIpbWkIiYSkDgn1eHsjXq5gpPvjq
nfYWh6JGObwqQVjpPV/wTuIOUVLGDq8B9Dm+25IYOZQgZPNeq+G5oIzjJbvT5ajEYYuz+1DI3EuI
UGuPNICi5478+hqW96rdqd+NNW+P6IPX0W5MW8d1M6CwCjsp+99b6BUYlg6Lb7cCwJ1SFW6Gcr+j
ReYiIUm5ddubooJPfmKxJk13FTaRhtZmTFHxFmGxhZo5pMZZw1JIbwc/o0NFoeBuXn25poGtFS6m
8x3yV2qoruQvrPq6lZlUVGzluQWR09QtOYZFxaJBU8+n4KLnE/Q2iVMfoZTyW00il1DCMB2n1pcE
uzJbR3bQoTRRw1IVrIQuZpH0h2tF21NciYhsH5w2UzH1ut0yMZ1oZfIst+KfXu9JAvoOfTBZ05fC
MFe5M9LXfD4g7qaM3x0OyhWMcQtGRiei0W1VaqOdA5sOr3RA+oCpjsUPE0Dy+fTQkt0cMdZmBTMn
NUE7ZoMS2m6P7UZNd6/E0xXCKlAKhNODWeXD5c0aBMH6Iz+3BGe3Xhx/XHN0N8YiXM+sPCG/diUk
FBe+jR3giWPaExtgo5pAcztCs+m2M9ayIZ5OXHDza249XnGoXgv3xNJipeaAqv5sUY3Nvkp9Yy2w
zUvYukw1QoKuaVyp30k54kEZM4EUpC87N4E9Pgl+WhyhmTd2CyIpIH7JfK9wfdT1mnH1AGBsssvb
cMBY7h0Dlzl2BHRdf4mUpuKcfCTUwsbYNWm/CYcyCxVoLHggIVNzhnSU/ZtkzuKO5PkPnVX3q/fq
FEau6yCd0Nzl/yVHKZR+3MYsh7bIGFpvQ7S1p03dIrxt7BepY9a3dGKv54LOFSlXSnnZcBIdMyYc
Phx/vUbK5Eyxpu37EcC1MN5jb/p+1LiNo1qmpynyMQa7x0KmQcioUzaN/4/OsIewmm8MjPWYwvCn
qigpyAZ3tmObLE7d/iTwEJ8RFDw21SnPbgXtStSekun2tpm/cgaLn01KJzeOxrQ0il5FXTWwqdVq
yDUxo06QR8kuKEHB1UIs29WVHpDG4EqgiSR79s7yKzpqg1NXiDFtKX1mTnO9McidXMC60+txTKnU
vSvLn8S5am4SMNJAbi3mSwvlHfd95OTllNMLO9rR0qQRzBBQntZLL3pBYFP/CU6jvGlDGLhlaTVA
ZZBe57eBICtZc8TdCfvvn+MJeWUNZHV3fvMqUrrtOrP6L0RonA7ZW6RRA67yYHTv7jFmlq7Viyd+
jAQHZLhmb2TxsHpicxLriTpOlWs08o1hxwCBiVNazI6GNrouofrV3NIyM16zGT3xCY3luV0ydg6m
LIJbcNMEslD70Jqcu00yQSFTusSw12O2eREmNCKL129zjEmBqstW3ND1r6/UYiQnXqMUj1R+qU5U
KY/wTuEzdFw91t8T3oN+rDeIx9NshEtlq47VslAUznCkWFm4tGh1d+C65t0nqqGfuuVKe3K7EB7l
pK/uuI1ZIaoCF1czfVbKlVitGdndSJ8OOGMeiqRCJkdVk9YFK6UXYm6iZaE4Zqc4lNsGjQzxWyNG
7maJyFvfWjoAy5aBGGhmkiUZaHuZsV0FRz8TcBbEeacdoO2drR8ZClgcYm2mvTP5NCx1fJjUFp9D
yy5QxVsS5bavwedeFE2su9LnJVkhf2ifeZvycwSEpwDf1KtEYevQfpecGSh4rO6g9PbzO6hsZn/0
zob2Cx3KssC33aL7vE8L72UsK+nERXMkrtU/xM5WCNM6RlOLz+P1lSiUHo6N3tF4S/Awf4ePin9Z
NmXfgMEJU1frKK9aKo2X+ZNwOx0ELEXHVLZA3aA/4A6QnsqwB/V+sxTvjayA64XYM4ZYCbfpZNCw
cyMtJpozzQ6RboYIgn0Rttr8V2eukTS6T3Zuga0inUe0zfv2Za27N/jZ327Wsv+62/g29thArNgq
2isFTY58BmkZxH5YaceLT98o+lVOEBRYqQG8Dgk9FUxtTbCcxpn/BcGyssgX7b+tjknBCO42AY1n
mhJw5KhdpN46g4g/Wak4Y9300TOJ6/h/+CiEA8eVWVYoie5gDay7e3WnGpqB7A3zJy8hmOWCKl5v
6PLk9Ee/FfWAX8RqPSdRlqMaxSneogPsnand/jQfMVtYiVn02T9wdQuDrsjbYtqJPNDPFe+jDwah
BlWuOWglDV2/DQ8+mr6CTMsDHWSPmhFE1NVvMvAklklKYz+6pML7xAsSjuru2dpqSyEWpVCg/q66
I8uW9c2jxgxJo7vG/9FNPdYKo00HwZgWKdIprqWoLGH95fzUZgRmyGv52MicJQ3G0eKGjNVRFJHm
HOITQM5Px3HTuKs/WHn0ZbJ0Fo3JfJNxTxYM2YjlCMviVnLAg8KdUHF4W00+YzXnoEnGPt+RiI2h
SUtDJjfFVDFQOFrg+ODGue3T9G4zfn1AdmRR7wiPKqCXmoq1zzjlx0WYggxoCVtiFckecA+AxOb2
AZw2hIXJigiknR/tuU/QHiu5eAQkrODx2XKeHDNYoBHsL9e2xgio8vYs6lsmeYaAQm7ld/tLk/WH
aYbWpMWhjCclmf2dKjbLCx23UG4ZcNStVRVlXnGdbrXyfNfGmPDgy5d5UXtm5EsiBexF4HA6y7ja
FzoxofDwFvieXqzkBDzTKg460QSYALI4OAFnH99Z9PSnVfhN+2rGtdTFe08xYjb7xYsqX0EmPaaz
Mg2nqafkNC3SZvI8AJUnUn16Mc/irsYSJlSjsXnvDvWoAKLYrlxE5Z+WRzCRrZ/bTJahvIuVCZs7
GEy/DGXoQ20SWiQ2ytRgYdJxUNyHNjKhr8jkVzpQh3DGJ4nDhCn+yXog4w+KEXHGEpoHrM2xGkSK
TOblh5jcKdiR1/k55cRp1KuVwV5mKZsGC6hPdhBtUzZ2cAPvZhvWXkDkWqQwLUTKtB179bJWd+u2
jE/QY+bXzqjKV8YvF8a4ojhlmUuNzPzsnpXNJGLy0Ccb+FSntrguCPFlGd05EKgT1eh9M83cRGtd
OiCzQaVlvprdTPtAs7DpXq2pV7eakspAJ6OFWd31xR/pmRpRbb27eNnNSs1YfTTs0qMyI4/4QyMZ
BupEVUudJx6lGuM6SFCSpwqc0vJUexXJuKyIMwZIqsmu6awBFM/jq0M+3ZejKRBo+jUL2GMY+/yL
qyckQQUzY6t2AIOWZYIaDKpbLFDbL3FRb64y2Rfvxx5Q54p9devBPxzh43IbhOewDZaU5RFiJ4Nz
YVcnBVu/7qovRQIwZNWfdoENVZvmItM/wjdNBL1tJy7cizD/9iSjtar5DJCg/bYEw8ACic4AnMmU
3I7kBaz4pV6PcmuXKwr5VYP6qZQqgWvetR6WO1IrYotruC3DpVfVWwtHXDtzF6J0MovFszeEATOX
SbgRDrvDLD8BV2Ouy4VdtttMr1g50c4f9CYz0I4UCRxz+AZgcHPQP7T2xfBYhwHbo0Yjmcm/xd7i
9b0RONDs/EXZHfdPF0FuDnGvdZDhtXyYB1oyL2ZJS8kNIF1+AmsfOU2310RKzQgegFXTbfvHA4+D
vIMK8g9xupWAwmu/Lsixulu++rdgXq/RbkV46oAm9oG7F/vBFroK5aBPCsVGZ4TAcK61I3CaJAer
xRvGMW/WYHhov9Z+bm8pW82A36gRFCB2wtqMZ3H1xYvKq8LeJw6yoawU8cALMyIM/tOT2qmiY5bt
3jaUpr09oj1mikonHI5QhcgrdnWoic13wgidVG/0qjPktaapoLrsAtusLkicY247sZId4K8Jr5Yu
se615S3tPtU+GJ9etdYMqDY0lxk/pSYCzWkwtu4QBngeflpG3khyd1k0fb+A2ZAxxzgmPmGfFSE7
/ROb9bHf4VzbYMhBJjiQUwtH29N7EXe4lQRLgzlNPcvzFY45xLp/gOOAx+muqGiiitGtgzJ1kSXy
88UnC/5iASSveUu7jPRMFPesbev7G2OAHn55SOXWPIZr0rNyfmNiJlhAL6htFhs6CkYpMPyD1xvZ
xriruaQuZtAQxbtmlcHwhiMzW+d2BVDDrrY+O9P/esROD39+YZQeLPH9gwHl+3oIrb+AuykfN5Wy
NCkGQEEHrV90AhpG43zBMBkb2DR+pVlkA7b4E7pAmVXc7FBNmFBhFUDQzRgMc5ALRzwULgsGIhoe
6dwxIGWRF/ri+0E8UzGypW1Lq+LeE3PQ8F4Q24fhW1IiLBnL/YemwExx+dWguvkqbFj+DiloE2CO
0d/x3i4inLfZLiwhlzQnoKs1TO2bjuX+O2oYxwp+coear7Lju/ihox1lYnrXwG1RorGoizCvtkjH
0g/equyvMqs+YmmhGECWQy7CsA96rM23sQn+9XlFV65uUVXHm74OX6m4/vJAxWLCIWayZMM6yTku
SLBYk9LQ/M3Ym+qyq1QVgHXtIylv66kjVIYHYrPJB7C8BElH3/LuMEtF7PEimk0aOCdQX6YMuofy
cbZl8x/AEPRQtKh9lBoQmAb1BYEm6Kyv+RnH+o4JcJezj5ust033ogVzafNn+pXS8DMJk1JTeOTH
BcSPF6DCiXaOqf6zYziGdAmymEM3E/lPGd2iWhlRc6B30NNKnIaDkgBODiAW+k9Tp4cRhla+Ghs6
zxEI4cCU9D3Eh2JmjJmOV/za02ESZxqMaEyPKe3yrK0bYSztMinDZ5y27WPOs9tzC49bqP+RIT6g
ewfUFvhEHi96VEi/jSnnO3Nm3vrXP1fVGxDvM50zBe1TtMzBaFRBb0MRh2EFuLmOpK/ZMT6F/peN
v8Fe0W+mLODBWPuolL+03hLOZcgA0Nx7I5yXNx52LZodGn03eCZkT/m57qazYyWnAF/ZQwy/aLDi
SLaFMVe/8kgGvTSGVY7D8orgcy3H78KZ4vOKjS/ysoOfNywJiQfMYCWBqQxIdu2YPQqMewm0N5nf
+13E/sRK7SCipmQ0Xb+pFTx2JjGpJ+DpIcaT32hTXfZ0EBWC+9noQ/gIN3wy2j8/E6xuCF/88yID
vZi2Hgq6lwDSYTYpuLUDXlpcYVqczB4Pl89jxZ5ikOi+4VOzaN9gqzQDVM2nLbPO0FWKZAzPS69o
ZTIIolTx+4Irpw8X7JCvx7hpX4yJ+zXWY4MscG9P23NQEevLJSHAiYt8j9qDW5e24tlkIH99oiNQ
bn4aOuixkIrp8p0X95NJqAU2RhA/xy2TWJr+L0bAVoa4uLNDreYfyCvYN751AgWbbvjpsYspr2hl
f30mHy2yb5vemXTFC1rNPLgBnSQRRciJ9Z+Cs7V5F57yo5/k2DqmWeQdL6g/PSO1iT5uwbnLkoJu
hftFPsqKl7RzGmohY9Uvh9oYP+sGSihu7phngslT5qCmRsStG3NX+TAtRv/W5XcGeIjW5HZ23W+0
kSWXlOD6H0QVMF+iNUwsTfLwk7NjN0Mxfiow7kyPVXsS9dnH3QxahXeHv2zPvURwLiAVio+fnkzN
DfciSEaUPVajwbnAKPrNiZAKVf9zsJ1qogSJRMjTkgh+yWGdp1uKDIjDJolcjGBQoA47AfdoEa6p
vQSJge9hYWKj9NZykQSNob4iwEXwJ0nJQTPpi22ZtMQMzmM4KgT1K0LPjVDqUqN+7KXEXMF9UAuW
ZgeZVIomu7XC6l3V+G0sGL68czdSIpr+o1lx1v/nQFiKD01vd2bqMoBJ0Hd4Dz8dgZSUNWW1+OUg
y4vwkFL/unjCFJfqf4Ro5GNDtO3hXe4lcHqdM+1czGq2GE6VQ17mAEqlGjfbvlwIAH2C47A5UMlU
Dd4jStfwHO3yDQcA04BDb+voGSrnX0b4wuGObtGY7q0YGRp0aL60mlHjFWzy51/C/QVrMLhZ6r3s
nWfW8D035QBmwJytNmx0o0KcPDzweZxoUHVUSslGr7RYuI/M6M5gRktNHZWmv5wMK6TtPNTJwHMr
NXSiXMOZlcUI5hItYitJEjktWs/skay+khbf/pMaI1zCwh7njbIfZnrZkwoCgaN476gbZYjhoYcu
07T1jYhUERPv/kWdv00/op2NY5325eqQfIuSRgITo8aD9dicT3eONvjE1mw9aY2W5ef0CUXKEhJo
A+rf9gdAGoyH68R/6Yr7C/nfiyo7q2G1BGetPQd4macDxouowTWflNEf5WiNVzOP7UnrgGIg0XbW
TbSaAYW07xVhxD/JfBlVrMBqPlj5wry8gzWQEpFcuI4d6HgO1yUp4WEqCRAnvOkjnoQrhHkVnTsz
KaXAJbGSJTre5OogOI/mC1l61iJreHaKSNee0VO6vmYqcPUkd465kcRynEjEFpXmu9HsuegqJTLa
M35bvjOJq8glarH+Mb9uqif/IvF3YXMz3p2vKc3+zVD2oggNvldndTnxZW3LKkM7W9NdODd7mgKs
eokqQoqT0vTGI8aZ6hli57ueTaZ3iG6Gs6IxdMM/7pbSN71qKtPfcOsxDcRnxshei3ce37jgQuBI
jBHQnZebb+ygiPGx25SWXkcFrX2e2SIR0j53XR+w0iod1h0a/xh3kYd+m6ZYEV65sx8mmXoniQoW
bjJjtVcrFcjNeZ9oRht5r0u+aRl6SaJ4pr8+J36TrHsodk74/jJ2j9SpAnpV6NK5O067V1CiwTQi
fZ8Q7hBnpjL2kONoY+uftMDznbGa4C2LXmWhcwlpocPnNALRKXk6spYevBPIpUb78aMtTLXA5iFF
eoFY71No6HMoKOQKpTNfCSvoM5A9KfdkOWmZ35K9Aot/WbB/6DEkeyF9VIeN4+ByyyGxkZ2L2Y61
U+WbhlfEsLbEfFFluc7VqFuH4+zVnjETLxTbnDrHSSgpdL4Cesef5ADADxvItcDoi0LIa2HSwiEa
EsRSbxtR3C6na5SjvlPQ6hCeglPP3+mF7MeVbMnpsIyUsliDjljBx+fhnSMZmpPofTcbhTeDknHy
TJ0pYdrg5XNMsnA2Cd02G8G8l1NogjeBsgL3YZtauZZaKYyDeMeZRNzh5pI64ahYiAiT4ErOLtNJ
qLuIEj9LfVCT3iJ4Yy4N/Dur1o5999KxzqMG9FpeqfCcoQERAW1phvF+/HQq75BIJat5CuyccTTs
O/nRq8+k4wGls3PsUVYQWHkx+OVbD71mMXEwnTJIf44pMeU4GhSJklLp6J7gYAIP8eEZ8TeychfQ
qf9/jIPxYpEDI2GMAsVsk24msMQ2pTwIvfwQBM+qHN02RCM2Um3HQWhwyEFzV1eeHN7oWjhaVsz0
o8nac5/R1ledJY8hEZ9AHVv07tWv9/1SRTEp52GpSJSGr8cmJKaHzM3yef0fZPDEBrGjTSN7Kbvy
gI1WwHjcV9BYmOzcIqSSO0uP3jkRSJMnnBKdSHLJLbwYqsVfgBNHVn7jpZwCYhjmJM367J+Muknp
HeWUhSvYTcIVoE8Kp849hho1cj1b9D+axAGQ7Ieh7peLG8a0LLpkTs8QQiUjOtFu47/8ZRZn5riS
WKggb9bqslZv2VZ5TVSaa3y5qhKWzzcqL3Xs8R/3aU/HjEZgucohAPlbdMyofLEhElSyX7spYGdG
8kLX6TZjB23bRnSOytBOytbwUsb13ey565BdEMZVPbUzKzCKOj8Y2h+qeC61ePQDh2mqHpHIpnm9
0V6eEpPX4gfM9ZkBpWDykEWI+/72NfB5QNlI4XkE8l0/RLKNoaTxP5ID86iT9WP39N/XIkGdzdBN
oZiHkR7VW0KRMuFiOFClc/Z7gb7LrTOG8d0Xr9FLIkGPwXOuXh2UlRMxlHxDVLUeragkPR+VeJOD
1ldn0ZSFL38DtYSll03/f9dIfFTdWEnmC1Us+VLyFOqq4fW1OKIUY+Uv8AoHOHf09Tz234/u9FKN
b4QzJOhv5G7aSQ3Qfzh0hQY88Q1TcPjBlWyTgAStYXGZeStUUXIXrcu7DwIs2NPlcXEuFuoB4eKO
q7AXst/89D+BS18Ol5CGI+pC3DpTN52o+H4/8dEfrBBGo2v9zq8R0C2FqZOXzvj3aDva3qxYjx9R
RY3COUMes6XkR9QwI3RAh1Ru+Qj39sRYQwXqlQqN/B87IW2BARcwE52MdvCLmqZ3SElsBQSDBxaX
6CI8N7/xMnXIHnSIYXc4l0UDy07yVTddslvDsNPpXGAWGPsRPncHjcA2v2BbU3tMgk6j1Hx0VHSS
sNgYqTRFmlUpXTXqtoXuIDFocrR2mKQMtFkWdX+7mdJYJK3HOyiGzt/5CEP79CY5XjavbAEutqyP
59qmBQpD07cV1oTbHGmDsnp0g8fCbUNOyryncMPNVOlVqmEN+i7q93DsLF5TUya47+A8DvFfPDuD
kkRVJfEn2QfzcrA+Ogy1gBXhoSSO2HwCGrN4KC2NJlq7GaIfVz20JQbts+0UzMDLyNG0lNCWUvtB
uwjkuiUobr+o5zPtl6PD2OSigDaHis6I+5A5u+yfJf36GlIxDDAkPI+8qp8LTvfTPLBDnrW1DVwF
PCnGvi1g0iTF6Zq9/qZWCqaMc/RdvkgBcVsn9/ASy+aQSyBI8XU0IVONgwFQsAJsZiKTh6cqghyM
sGv5FLIL0pw5wCia9k5PcTTtbuRKOVIQ63OKC7307M93RjYQBM7nMDOCVnT/tFVAAhOyBXwU/Exi
2jpfS9MtsGb726OKBbdqQatI4yImbuq36B08JQ73ZBBV41rWNPPmf+Lu52lsmqIIzPny6G2YKVlh
QT95MCcapiqhlDRKzwvDFv4D717pFfto4hJ9cDMJ+uAZS1ZQoAX4+chupxkKvPYriIQTzI+TWKAk
RGtjnswHjs8XJdshC57ZO+Dj8TOZCJFBxfpMSBxHeDmcFDRfiF9CFoXSEXdLuTfyujGBZD7TCgUi
wgXuaOvJACvKD4cmXwbKyKPqcAhAkdB+xJBs+QETPSNGs40LIRiuVJkVEVKHaf2tMPYQP/JE/ZYb
qykxDSpjYzkvxUqSmEat4T7pssBA9LbhoQyp718aLrhPQTfxY/5vEJM5tNsPdrugwsGxRzMaCJmp
dnlXN4RxJV9HXiQL8drtkm21fO/whHfDv0WRg38H5Cez1tVaZenrCTx2Jx2TOyy15MTFdTdAOfPw
Qy103EeBmOD2v63bI2MgCa1/XwFcHF3wVNNQ/p4j60HSs7cfG1/h5Wt7fZWY4uKDY2nZmyKAGYOI
RzoRIDALXqXVuQWNtOomG4189MknvurPK97AXc47UJ0z+K3/WwHFdyBqstmCgNOiqiH86ui0UINY
g1SGXma7ly/w5DLr1/Mdx9LDusn5x/OOMIkQWt+kFoetbqv+Zura77SopUx7JgWJwqU0rORpQ65q
0zE4dvxn+U4cGKzZWxFxmO2MLQjoTvNfSfl1DVlyGUlDi9dWD3V7muNJMx5uByxLByENaV5+rkH7
AXqAboPdcXPD8VvFTH8S3tp/xW3lYlG6ncznV+euIe6ANjKqKuq8ZBw8km//L4d98Oah2D/zyN6z
I1SkJl1EzEg6VrAzRjqap0lKV2KYP8btL0t0+Ee75hIVBW0MTeXqxWLku1YaVTGGDcBKvXbXUSY7
20xjAyUh1BZwrgO/Fwe5Oky5IBek5BegSkfn4D1GhZoP9LegLqLSeyPY9+5klJhn4tLjtjqhTrn7
6Pwsitcg9bS1FLtLdI+oNkPnmD6NkgUSsm5W6Nir5D7H72FE3d1Dp0/kjwDTcuZ9nztTS1l9vQVK
phAuTbxKJg3aLbdWbgFVQho4gmyJAxERfo8UNV798mQCZeZh4xJvuO/2c584J3bey3bwJzz4l+Hr
AIKmE55grhpnynN5AKN2oaDjlrHVIx7TFgrzr/StNJpPIvKea28id4vKM5BNTgs6cPF6ovL5hWhG
s94/1fIq46YRmNbG0bYMZirYoEcbELFcDE9y27WEsxQWWQyd04NvgCcx1CvN2nLSd9twhthbYAK3
sF+vn1YyQ+TfREg1Pi3GDIdTlhhM7tTS7Vgqd6O3dGHlHOCj7wlfTq3GBNzKucLIH7SyQvWbiH96
p/q2kEbJsJiwvXhgVkBdv1F5I+ZfMzKOKfwcpGQSJ6XXDMhbT2WDyTOH2pJle0FYqtwQEUQv6Pri
X+UF1drJ5rFdbmOzatBCKlC8x72j7cYuObm4vb1BjxiKmMUbdHfXUmwDFY2tppo0qqeX2jTlItTb
RYKeaZPSwGNHNXDASE62t9wSVtXB/T5Tbg5RhW23ZunEd88mczI1tII847ojRefb65i4QaP5jAjD
Mu20/fBazQwcNPCHowVXUrGdpvd/26rTeFcwDBGivmbEvw+tiUDczLA37qAaYjx3p1cDu/Mx0PEe
/C+K2974JNxDgPPaYCVAWDAw30dr+aUcQjTdkEqeinyvSyb2XYlJYIvKezpZ1OXAXE8Q6ppdHv21
HyXUCwNWWD2s+HzbfCBQHwbHTgsS//Gfv9rUIWZELmszV+4B5urmpL99edTPnEl07g+sw6hHTowA
YNsG1zgfdMyvR5xKx2lgQ/21Z3YkPCyknNs07aneGbu2shdq6oeTy1pTwPzYM+E90HVgXMvLXMuM
ud+OIaQ3BRCxC8FFLZRviaQV2u56muloh5gg0ybYaGpsPTH/Llb5Vj2Uvi5Jxs8cGEBo6FXuX6dq
9+3zwpOOnK+8/X368ECcNECpXst59EeRxqWcsbgU8wLp63YsAuosZ5VbTdO3OxDJ1QqOdYoPkYOk
MtBI5U8xrgFmKCubgpdg3zgK8RBl1emgbrX5/c1SGsCEOQ3EX95X5GN+hD7icofvdVN9H8PyjAtB
MqYgmYLGYqbpihV6xjNR1gymcXlW5VzFhUKbnn74XkK9mV5QVUJyMKpPplZiW/hww0gnlHR/tpaR
7mf/eBvlFkyviWHAhK1pN5XEh5dToxb41v4BMT/cLQm3f6A6IpORMyOlIJURyfPlbWIW8Kdy3bny
QBNG4qX6DePOivWVU6DRjWeuhr2M9nX+0AMTgy+AW8kEjrEuQ78LQzjOaZWbUnXw1ZeJLW+m3UCY
OHstVIYgyoT5UU51yf8Lh+E88/ULMzlodlXxN5V/nqaUM31dXpRBlgGbyYLZQAvtFop4CJmj2TP2
9+whWwJYLACW5zn4HuoR3wGG8NS5xEkjVXTHOqArVy9G2pXknZPmBIghn5WUcQ9zaThJzuUylSx/
aleaSWDkznXN3kBEFBLA3iJ4kxGKOd/3VlJ5m0MautRHtKWfPK/8HGE4V3dN2Up2Fs35IVFR+4dG
A1mPf89I+Axm5SW7oQj9TN5AS8I/h936xsPxboHQQ2/Rf1o0HZtHphFi8qS6QZ1QckxRD20MAvYX
xPNbZJOHE0p9VNmHXB6VJq0WbHD0Xz9RaV4nB9j36KpUbW/x44XG7vR3m1QtFUeH3gyHI/pl6FDo
faPzt9ZMhDR3JCbSQRPo79ghSY46dtadGSwHDhK21EzqOHTVjjFhIaQ94l+gF4E6HktkxqRklWgt
eustnD2BV5+Bx4ZZyyuQxkIACSomToyP1cVVGEdgtTiMcRNGAY32YBWIfWzLk7OrXD6NHbGFpi53
jLkFsi38tzIhsiHbcC2UUrAmjf1CB5+ONHQTe20VT5W/HI3xoq9cTFOF4C/BvG5QLyGyEhiPRxlI
1DIk1kpaXs2vj7nTWaykoxuyqqB7DG3qo/rHhkYR4mBDCfN4HmhDV8dUVhRVhz/OlztCPZ492Twi
fw2z+qUa6oxrP8tViDh1bE+CHsSmb8pBfo4h402MuC+PQrlp6oFLGcu3l29xqHp/IGeNJ9Q5PFPd
f62JqOubmVRg3sUoMI1IcdLthj8brJOLXZcC5qFN8Ttnx6EZrtDKpzRhiRkqIudvqYOKYrhPQdzJ
N2ksrUXJ82kOhwtSQsqcSjG70XWD2VKTraaIsBzDtRCstfPuVEVSFI5262ovIFA+6q9Gd/iHiofk
wmp78Iih4moPue6BWRBnBTXY3+VTe99XTUfDUTOXKjoOUYFuP9QK3rqGkcren4YZ0sndExakQDIb
XLy+zbCvr8NeOtWSCbF67v8VwOUlyI9/EJXKq4OK2iGoRfQgZk37sT6FYOWQ4bmiLhYu+12ucBXx
kZKQA1J/iTPU9uCW5HlEAahpEQSlQCsnOsSb/iDahfuUGh7op7dHMF5JozzygR6nnrzAvki+WziC
wvMiXAlTdEliUFRmR062MK7HiM73/mIumeZ9pDWKMTt6LzJ21zo9pgqEc2BL1LjcYK/z0phO4Dss
5SxGU/B3jeE6zzlbztDqr29qGEqYNzAO3kw7ueBOgmlpFDTrtG1CYL3vaYHfj5ePkv1XZLBGXsb8
x0qtHMhHvVaoZgZMZ39EcHkAGnSiTThtsNx73okVN7GuIk6mh4Yq7YajFiSP8DxAaLuyEjkrZDPo
pk7WvuBRxqtTIL3kpX5wJFiMkHa6SleBcZurb+ECV5ocAUJJ4DgpBkgrZA4Jw4Gq+Yeg0/xuCHH1
OMmcd7QHr5C6sEw7/3ZlJ53CAClBBYH46vW4BTq6Em3RWKu3QGKhAuCKVkjyNA6fAl5Je5dB//be
BfUUmXdvh64hfiCVroy0gKGMTsLnaJ4zNtW5ygi9uGwcOwuBS97X9ZxXiBgb3GrpgjILFDSfx1zA
x2l21Wdkkmvp91t+NPdZ+24O/oTssfeTU3DbtIsOuDod8v4utj4U6nrF4UorRNwms9iohmv9rDo5
uLcAwwdsP8EANNmX9OaGNUXRjTzkSBLhJX2geJ1LbV9ZTAMRQqTfBtedsI1QUww8DgEiKUHZnF7x
rcaS2kns7KrU7rzh5qAajJErRGb/ZhALPKnVyBW6oITGNLuFKBbFnVjLozYmPNKapQwVpn4mRReC
uCequS0igNwawa8W/qGZ56gk43gZ+g6nINXJBpKfD6bX9iaR9RdBhGXuVvYf9Czyxmc/pKIsqIaR
8eCzlzRZLYZI4BJyOtgOR6qsaucdOiXFsOYwYZclZTJU4AwjaQDpkaKS6MkEsv8nP5WfiWk9swSq
UpKXbyEVBOy32zQ0rA/wdIpkuViUbueSIsN8YbMbgqAwX9uIBFSbjunlMEETZ4VsHIgIHBM2OA4L
4turqnm5zcsjdGT67ItXHXTHezGKGDwhOw+WIfyJ7ZUdodpKwu/Js9U5kjSz1jKL7dHotEuIxitZ
o3u7K3DVVB8wKqIpr28j/DNvyIVGO+rQ80VEdMfMYfVukp1RY3We+zs1OMI0jDOG64lwxeZEyzZc
CJ4+VHKxcMp2V0eZCdw6jjAoFiO4FhP/1zDdikPw4W2fMjRSvBcmDzVnqDKNhSQxvlDT2Q890Ik6
pctgNJNLj9ASxj7qYbyIqWRMa78+wWpP4oGAdcJuIQ2Twyf7tNoEwT90M5k25yMHl91jRgfpxW6k
Dbjb4kFDhu0gKc8Vk9W+OPURNDLEWOIfPbEiiacDJWa9Y0ivNcI9N8dY8ZrWPoJuN25+2bgVaN+b
PNLR8+Zt5fr83lQl6LuuA3ZhaywgqSYMfpdNq8inFh2CCyIn+OuUu9MfUxkqE4xQw+meYEgUp0Ss
5ljVBe24VwgmM3J+/lkHs+YyOoEYExpm85jELK1P4qSyRAfXrOLC60R4+9+BOcNf9t7vR5FYKxnC
ILtGsUsGBQY+rggKiq4q12yu4ggocgKtNiotFJLGn8t84j6Qt/9oBWaz5vyQaPzFBV7oE8Cm7mUt
3ro5dCXs0p5/WSwcaYNBTu3IcZYLfclNsXNnJs3TmDO7L7jBzJeS2zdMoYyfhlU5zkLtc3T3s/Iu
hnHWwnZwu3iHaj/KqnyKikUP3mRY10DHdiAdw1N7gdmgmHILB/ejPZjIWEbNgn0rm8RH4NDXRAU7
IUI8N+3vZWZ6cjf2OvyLBfMXLGbf+B89WmXRLqtecdXkGkE2xF0H4/ws4/9a/VCYRJdySrcIlMK9
b7mwSPqUHbXu4V6zG+5K+Py6q11h+OB3Gi7BDcegxUZ1F89xnsUjx3fJUC/Hb4Xkm8N46jUCHRyF
zOtbu3w5YyU1V4MQ11iKMKSImxDDFMxnGyFOF68gY65nxsBY2lcAr2muVOZgTwqH4Jr+1EM+XpV+
h6bIUG6avAoaZ9phmma0t2aJyRgCEOGx5qglW0ou17e0ReDkBAPyK+8pOvTpfpe2sNunXNF8cryi
yYcLNsb/7tpT6XlWjr6EUwlPLMnTIanzQ5dSTyFmP+1I7BgW7iwCmLtoCrSNackmxpEbKQRDnegK
5Ujrz9jlKINCMEcy+Y+mMeJr84DPPYu4T3x23RFxwLvE1ixtY+pmdAm5zuIHhGrTuiPrquDEDffQ
Lpv7BAUmIL+vc8dkS0YXr0S9tllUpPTHdDQbv8IvifGLaegSWOOBQR/reTD9qRqJFtb5RibRroDi
EFVCyceb4KK/5rToQtuBFLZIF1Z2eT15xWfMpE+dI0cBx0u0ZWBqikKSlLdBHaH1OsCjSToHd4ke
HLetd5/2hKZq1sE61ceIa/kyvVwlS7U7VRBQntQ60H0Lz7zC/UCYz13Udp14EwyiwZvAc9t/tO/e
t3Np2tkmh9EFIVXGM7T9OvDJ3ys0InybGE6x912tKaOKvZmL0kfehAi8w1lAyzqC3Gdr1RhecW2K
+OSr8t4GCRuDvyG0NPvqsNG+h0fRhfQxAXJ60BD69m37p5JFvMXbRwEPLOrEk79Bx1V01KZC1HuV
oG7a7rhd8tfmakiEECfMRwWicwHRnJM2x5NrVzmknytfM4b/JHtsKsPCubODNuCq0/JEphP1SUvB
xXZCndQu+cwWE+F4WRuIYuj8LeBI3e6nyWmH9Pa3aCszmqbdE20Nz8j+lyF65u5SxQosFjU8i1Zg
CWbtQskJ3VEAeACiggfG9OvQ1P32jI3QjBqTT4qKzn+Y+vzyTNnmOUH5jYEjB8rGpU8QkD7BuNPx
dxPGpTgEkWW7SP6N3yyOp0aLRrU41sNG9o5x/1Q/prevrBO1w5Fc/7BmEGeofStR/yY/dYGPUJ3m
FsXddt1fXRkw3HAVotUV8Reupjyqui1ZVhvAM8lbuvaVWjqJiULbSjwu13EugMNF7hrgygXUTxz6
vwdOvGHce3NIYuW6x/N7TocvL0VQPWPMgj8ijZmxiMENNVG6cwTb31DGiyqJQ1Ft+CrlXAN5Jh/G
zG8dbwiE75xJZP+a9v56IelGR00VwZNvvpwP7n8GLcaYJwSnn4d5kbVF1oyyQC/xBBr23hnn+Tg/
YZ8vOjCQtT/peeJnaipmMGz02tK86eDCI+Ri3Nm+HFDrNr8D+YOaPza3N3eJNEscSg4Hxaw2IFHf
A29N2xnub1moRWOqNHXrnjwOmN6TyS9/8m8sR3CZ44/WkeIA0/M/9cxCF3vU7AavFsWVvhC2KUQ0
rb+Q1PKMCaLtzHyicS+EB1RenryFIEUyBF7NSRm6su4vevbwLoTrqSyvzgYoz1Y+YpzQIiSl2cZN
voQ9Mdfq9g73BuOZziCTc44ZMfzf5XfxAbM/nDssgYYSZX26jNboTynVbmR3AtnZP1UDLM49b52M
PJevUJPrltQMej+twZGbRbOmLH9IIB1XUNUJjGomda0lQPxvKzu/fW7drlMXOE8l1F1CybDe5w0X
+mTl1sXGArykCL6xRXG/1ZX0xqn1+CECKjDuGk87iBTccOR4jb48PxG2rnn2WTQ+1bN64PWvzePr
G73dBc78c8RyEgwbH0QlaUb5NJo+1X8Dh0M1ngd7nmUyG6FIStowWC2qtPeIQ+g/9nZ8xE32JUCo
EGp4h+hhCm1CvYHTVzm9je6tJh2MlIYg6aCsrNh4tLrSu3XpxP9ESRMnBn9mqQtArpx66VzXplXZ
j5N1omb7FQrQAKR6vfgqXOENnytk0EzZ3PFavG6dexbGKEJLhkPH6Dtl850o/0QZ8AfhKX3cKtDX
AHpjQlJivq2rUMqG24rpeeMSPnTiix/xkJbRck2rl2I1/qsKpj7tOKcC6aRPw0510YIL/K8ja9D8
du3Qj+lWNQAV5MjE2aeq8/Pv68sj7OxcQG50LI5iIjrWwu4Z3UFPje8Gs4QB5UFvNECpGFgI+wZi
mwzl7QXWhog3hWnxNJjxfO6TrjRFRFs5h+MBohFSLrFHzKYGs7Y1MxEkyM+G60Xi4ZtBCZrtutSf
xgM0cw1adQuPZPINoQJKt9A0hEhQO+/2TrvOdblzAxtSe9LQPIp6qYIPuEss3U7cx1DpBOqsMI7e
2WBBGSrGoY96W/qEefvy9WlvBF19RC0v213DDDtdo1rKJwiU2MAk3ep0h226Ks4Hdam9rOc/nA+/
AfBzsBnJr1PTL0QQoT4wInWtFkYgnc/wa7mELrHGHTZv4Jklti57ynsTLgxTOumr5K0TDvSXjMxx
5JTJHPUFdjTyBAcb49/UPfSnE9WdUS/yCsCARdnZ0nJ0gx4Zi+Ex6XUAbSDlNRgF/X7O+AWtOm2U
ecK2isjJ9+/LCIJfmN8iuFMOHz4/S3+CjJljMAT1APm3nj391gxitohLlY6lOkTgdmXfLCGxKv8W
2u9+TyPEDNRMUhr3ZWVsEZ5NiZDk6ATty7xIfjL2E8Caij0shgj1hE9JDGKA8deaf+rsBskX4kmn
ExumyKJJfbFgy6bc1ao8nMkxb62fyLDtYVyPNdp1zH0ez3rDxgZN450cOp/cwaaE5IndD+A9Ytzt
lE8TLPasigFDmB/CwQWZuhfA1mJyzE3dPh8IFfKr31NgRxKKvm+8kIfSp48tIwaBOYtvsOEiua5K
4Yv2kyoX87TBvsuUoeeQWKOGAANfYKKQFMSpQFKcBUFGEhzeZxnRFj/HGS7WUD8aQSnS1fpCFb14
mO7w0fk7MzMAv2UsPc9rmiJSoXM/nSN5YOIBfqO3NArXiDqV8DoWnFF8GHyhHtW+sZ9hYsqf0dRh
8qYyVTwd82BnB/niYOOQhtq7JOIE2PmYcSBjt+bHf9EnF76X0Ncx3ytGrxAk0xNHToQ7CzOK/hBU
kI666zcZxRaZcKPV6HqMh/m/hIwMyq07ZQ7fQfyJBxYkc2sWonF3aONeME4Ih1X/2GliW1N02Coe
DoqXfg/uph5aVYKLfNw0O97YbxtREbIGta5JOaRAXAfogKgGVO3Weqa3w2vgWIu1pc5N8Kgr2Ffr
Av1h+v443/yeZAPiI/3KC/oIR0RhCcsAuVbSRRf2Ui6n+g1HcHa2Y6HFiiO6PjxmfSgatiocCrOp
IXQcPFKmQ32gyssJ2K5QZvhgiejPmPJnUnoyoQRRclCS3TueeTrpRRdRUElALXln5ZFWKYvWQU9U
vxTruTeBHYb5cP4IOMFcGmJQJ1IRVPpqkdNQ6xwYipUsbZ9A1yvTnui72VfOxeZNBP1u9BxvK5Mk
70+gAZGKma4IDwPkQrlE9SFztg4cVCNcAFf56izint5dFuZ0xJAlCofFEdCDMsovau5glhOMjhpK
BsqGo1cQ3/9r2IDo9q011L3/nvYNqNUVyPN4U2ekZRgCeycY48sJakfq8cufGPyc9u8mTQ5K5KRp
SuTDHAfjvCh2fWyB/qeu6zNC5ZRXbtmIGDlqbyoYgLBOOI0303ruTjjlc5YKms1QBSmb4nzTvJB/
IfVou0miHRUhN4PT6L6ZoNfE9EdsMAvoSfZdO3uJAnP7bacaTICBLtrPmgHg2Eg6RdQxglr6uOHk
AZsgaf89w3mz+Vrp8ChVIdIAcxe/+KEI/Bhs74IkFdgzWfOjgdV17JRb/7IpYpA9Gcllid2/qWuX
3D6rjmXEFx4HXkHioVvpYtpzWkHczeCuRJN8ySpEiw2PhQSHCVDCb2DH5mn6i7kfFHm7SOivulpX
k8Lm67jBeBqVtXZLHprCiS25roBFyA8Jt2wyGN6JxVoYdSmITzrh0LSjnZxPz6NA/aAd0mwO4mEQ
vvkEqj+MBZWOL/uNH3GoTm2tBDly5HU57KNEfIfm6gjYxapUsYcfJJ/ouCpkvESgOP3V60vqBnQK
VNXFcvhnPutxi0vpVe9fV9vxNbf0PMEtzeYBDKR1vtiApj/KktJhFgXs+fyzin1Z7LC5bQF/TJV1
+2nHvBY+hCGOyD6I8LTe4ooygBSZ65KgazQq3pRKSQtSCDiAmPrrb/CWlktfBuhg7mb26HdTBXfY
adeZOhZZRn+zcp3xCtbqnyhZY70DTKV10wvAi6Z8kA+dUFx/bW3fDRqVstD77KJNcnUyM0+dmT1B
bW9iRIxP9dUf1PSyenRgD5CFtmCpvlUr8wWC+WpwOUCQ0qaOzvQw36Vj9vhAeqhAT8eLQth2Wiyh
ieDay8rdc+kF8HIw8RH2T4oeyNCIMCa2qGXu9uo3PIrEIbMbQSGidotgtiQdsvgQrnW+l+2m85Ju
eS1uhAuFaxkpflIhH9CJMpc9SIGW1xqDU9DXapMl6QeWidaUOPHdBxs9L5K6RGv1lcyJ0j5DyjtT
SDykeIXiFZzczhBigHzWG2zs/jE4plrTMW0Oro43u8kgV3lK4inX28JOnky7yBUfGPQArLY8xqKv
qVxyu7t5kttNKPzSNJ2H6AWdycTUA90K1W+nTb+1qcpiK7zBUeQ8PKLlTxYDN1H4YfWD/n+G9ZfI
u++quGkAQrTSYEHOJBOnUtw6QpMTZ3cPfYjkVUfz240ufG7ihWY47tX1bhiZWMUVU4Z1OZ9HJpGQ
yLq3N6bo+E5SU8aC0o0OagfeVpmdLPNktub5/z+tRzEJ2oNfxks5Bbv+85M+qWJ0RypidmcPeJs6
WioMYmoXQ7qvw+ajECgW15pER1O6h42E/MdTgs891sFuyDFcKKq6i49iLXs38VRBFoLFpHI/f93O
53xnrF8BATPEv3UZEK3RZlNSMnhPDEQJnHINK62PNkNSYPvp88pLArQttNMgE+6rWOnPVIk6BDiA
e6+GUzLE5yPDlD5ihCG6Q4TvvPk7i4Lbes2WcgJ+DAXyoSWMVUkiyz25os4v7sHHIMndwZHEftV6
FnrZty+MRf6WaIpGQytBpKS4HyMvgktWbwl9zleJdxWqQbbjfrRH7cMAHbLO+L9LOVGbLJEWVXBm
7P58RXXafbGeKl9u77dL3UuKDbC+SkzrXDdK+sx09DvzWDOJsJ4J4K9XAlAwFolE8d1bECXUqnts
lY9QbvWCFsGSZpfcUNHni8XTqbjc1sh9K9+/WNFX+9ii9EpDRVcvqhOvdBcAZEszf+oTxvlPnhST
Ae6FpOPCrLYaBayGO2iHNrXTLtu7qjZDw8vpcpxzFH00T86SaWUUe5XQgGeN4s4vWOS4u7mzQQ58
F9cVirRExtBRDlaiQpNAAY5qQNb5X8jVUiAlWWFjXy9V+IdivL5iE2ujEd0F+I8gQ5uJSbIBzz79
ywaiMvElgHpVG9L07vn2XWmIbrbcl8wzsbWkQWtqxNbwmhwxT2u+Q/Rd+dpE1UADc5UGREp6zUBk
sTrM7W8ksoBGt6IiAkLAt12BjFGVVqibpREKsqZBm1huAiEXvuNisIILjW565D8gptF/TyoTG0w5
+ebr7REGwu5Ho9fHHUIsNxw28qP72fd5jbw74Vr6TdtuZ/AaxIqNbKXPIbl885ZYxtCp2nVVb41B
s2tvnl3blDj5TzLxz36xjMOcvTIJKkN4PQvw8B3tQwTv9dL4ALSWTqcr0LGmiz3e+ed8dqDmMjPY
D+DwOgbWyz+NFHAUmhWtG1rGjac2MqH3+ET2rSOZSV7a5EKm2AIB8pH3NQAZ/fQn+JrRVf2NFLWJ
xht6cphSp1m7s6n5VsRK2XiAw3v1RRL4GvSw6tHfxlyCfw3WNdJdLAhYu6ZqXPhd/6n+VNHCscBd
DESp94E4k4GzMIxLTgswg5B4eng5zDN5LRA3Y9rFcHhzmswK9qjdKkNGrstIremkHo2pcl9BwbQJ
VZKpZjbkTHj7vmSPe2/QL/g7KeaaxQwedXX1AlF+A3RCSdTiQPWJyVyT1XGx0iJqaVqll4E9yHiG
SONarsEgKhQOKvENhp9b970tU+sy3DVgJShjG6Xq885Jv1abM18nFr3ViVa9lljW6nDYgqpUeR/I
W+YHJmySSiQQ0Sq8XtIqD/LSgAS/ePoEMunTOMejJtTKvE51b8nREpH3OTLIuIDyj2DdxAcroimJ
GkubkeGdePBrhg1jJCiuzVUf6Yc32v9Q/uE5Yr5S5KmmuFlHKzojiuAEPp/rm1v1mfyeQfZWfNFy
KONGy0c228xOqLJ2n/UjgNAkZSvX1J2h72wntiwubBnc+ZKQ3ZqWoWvXutLtzPgLlF7UDi6csYhv
Pk1kOX2QUilKp9lSxNmK4jSZs9dx/xCy8txBF6giZTRmj0QNq6Nsbp6mzJ5kKNYy4GXRC5Y7KqJG
Czqy2vBVhAm+0981u/G19CI1x4GBJriqc0qstDG0MYdvakuf1zQ4HDaFD7OsXFLmQM7j65dna4QY
+w+3zcbDztozd2hgQ2qsBYNQjMajClDEOn2JzfsqbuvqYpTE76ObpoRTlg0CPD04JpRQM0+hBgeQ
86gt1/GhWPwIp/i/NCt+vGZRF5/lp5Gw/IPKlSqjcGDELZ9AXuu67DgIUYxmSADx3z7jXSVlX9hZ
8c89+SrrBqbu6hf64ubIbd++c50tDTlQlfpjq7dy7iNLBhi/h5LxU+D9K6xUh2q1Z1epkeLdRV5e
dWfPKEYqcOR+k4sq2NH4vLYfKUt3ornHdXapXF9EOfHqSN9RNvGiDeka60pfF95WfDFktq8Wj4Tz
FFn1L9OBG1u3mVb/o+gd7btffi6Ut9zt5rC8jwsPodYpo3d2eTKCGPqs2t+E9T1nUsVRvZXPhcx1
nVRcPVbdXXn8+rBxBvn4G30fsuXOGMnf3Eo/0+ZKD4K6GwJrDnADr32y4PeX4w4ftOFzJb6OTNKh
ZqImCFymdQgJrGW2Eq12K+Qa3hhwqp7d72Rqut3fcRRIk3NDh4Euib+Flt1o5QKnXLlsWA3/RahE
QZQoUFAaxdHkjkCCchJID5/FX/QyeEnOaidVyq7RW33skGuo00a+KQCfzXwgoURb3S8+00xgk+NZ
IJb39I3Zf/7fSw8KZR11Dc3OjQuLuPektfQjZdXzu7eIIs0lk4rnBfktlNa7TOdtkrogva5+MjDo
HQtrNpETXGKoPFV9DJ7stvCpQ4Z6eD8ljBF6pzEdZFNbiqmqGRnZ+YPxIVqIa9INGo7Xhp77KhzO
g8qZm4YiIM4zTjUlfMjiCW+jjyk75iVC39+91vyeQNUQy35HJ7gOxCC/04LLnaWAhxYWAiKPjyoC
vg0jqn/R3niRor7DzUNGI/kP8zi/SvqspII/2tIu8+Ah1xl417dsfn/hMHW81CYjkLdgBtEaIDim
8sa9eyBEqmoNK5MdyQ2yuNpHbK31QvxAqBzlPH+kEFl6cmq9k1P2UfqGxNNb6KN3728K0/KLHbWL
ooXWLLYun5kBiwYxQszziLk3JOZYIAEj5zNTVQbX8SrTANy2YQjk+J8jbanudsoWaNH+g8/LOKKR
hmS1oqeI/696XayawACmG4O/G6yfUZGPSEScUa56hYns0R7AYFpGGr8jEoF09zxC3ZhcrUVZb2pq
mjxeboxzw9ZQAWFTZ0349FchNjZP+StvSVwuzBKA8bd83Q9rEoeGilpJBhxugQB38yGc803RMCFZ
g0JSfVyg3CuUlun19TXsoOQ27ZdRFd0Z3LRdIF49Z7kliglHBqZA8sN5VVEOvcldjJWh10f2RYdM
KQibCEYSJ/E/MsgCKxIFomYZ882JWErkq2iyB4GUXdr3C0/KL5lRPbmcctLyAduW8pXlCq1/mxt0
W/FfZx3/7K6/8Lxm4bc9n+zJKbZFUvbb9Ls6e16QaS2zRiyqrwY9TIXGeoBwcTczkZNxo0pTJANE
1Yym7PI47IklDVwiV6KkkhZBvKXI5T4hpJNtZGQCXNFOWGZguy6mFrnfCEuc/JOyzSh6s6JRwfjs
5jInAQ+V19N1TgemCrgngPvpuXwD8GmiNecluOawmKaM5/NfFUa20wnhwr4VnNcFVG6PVfqstpL4
Ef0vDZzPTsjmucfI3j7Ltr7mzCImdTiPokIa6L+FgBLeSeIuRXZLuKDvV5pugnPMOEx63S/KaZkh
Gi8ZhmF1XMktNneMD+UmmOfWvgDeo0xAoC6SMD9ocflFYU4H0kSXYLX2mH6JlSf5Ek1ZvicU9WGS
xsShqdFWwcEjtuKoNudCIiwnDKOwncgQoGpgoHD8JzrSpOQIHNyI7Grr0tEpxS+DEqTdROI0PmPW
y9776USs8Xa86BEesFGr74icYchhyCphFAOm/vULwi8+f4sDY8r46vgel3QtEJ7s+QmH9pkfmRF6
AdqPvmFInhWlRGXsKjJUUfPUy2BoxbBdM4Bc3f3+9bOZtzWSm+TL8nVtk4vVMtNdUUQK9nqSjZpx
OEI9EUuTYzdG0T3xMziVXHPPfLNCRUCFkMUbfcbFLoiCiZOwlo4RWOEa94MRguQx2+ifNa/EfAwz
LUzlxjIfFNvXw8f/+tYMu+8O8IOlw19CjWWRExzAoBij7/WfBE14papoxP3sZjp4rX7OOOa1pzaS
3b3VMyMQmMoU3eqL55gmmnVlXaSJzyGA/gz1IPCB4tCbJKSTSYPQW7YK34BFaMN6liRVZKY8KrTp
jguUbFEuOLEpC8Hiaimo4vFekzh/MySkQ0f2cWEo12SmL6YIAS2H+TVwDjcdO/3TXDWmSpauhFOb
M6RmauPh48TMXr5dOVfQv+8+DXaCp5cJE8qzpjSFMhvKT+X8C08I+mwP+fjo4a5RDeYq5UBiX70W
YbpEh7ohQZrQ8naFaS9tAk93iuxiVLpB8dQkmJK5H2Aifx6nQJAO13SrA190NF8Dh7CsrfVhAE5c
r501fZ83ybX5QFzJJrsZKmNmxOMV1ou0wHx/AQqqUoqj/UMcLrOTFn3coL1pUryModxKFlR3d581
Yz907557Kw6gvNGlCCYC2gExITZatU35XL8Ddt+LIY4A6Yr/MEOc0bcA3DL5srwd9JPRlU5hacSv
8gztdgn1yF3kBOLw8MqFM9jYYtvSrSKSqbEBpsU432QilKLnq3F5vR2kyAjpw7dnsUi0fjQ/K0mr
8UeNPWfBChIaIg6v12+GOY5A8AvmlJCEriZw+gdcqLzU/e/73kI1KufE1VKud2O88iw2tAdcd1zj
1LM0Jvw/qbtb+VIPT6WX31bhIXaybHwrjQtyvH6VF4pffqkz9F2O9EBqFUpwDAgj02sOn2KNsm7Y
0TrWrgbNGLhwIx5+dnwa6vHSOSSqMeX0mHnTxasWhs1G8kJ2Ybgj6m/TdTtwlt16xv8ohAgJQ5ty
b2vGKjavBKSqr7sqBQx2GM9Ma+yvji0vr6+M2iMQ/dzMBmEUnqu4OgtB2KXz0JQHQWdKQw2OhKEl
Ro9/mLimS1mlh9H+KJVJTXMNi2t8nHFf1iS2KtQ8otYozDtt5ec+2t8SqDEmnNYyBfvZld1DXgpi
S5gMk5njJSyqAJixarKHmAXZSAvsGlz1prMOkCC9V8PqpFNzckuDLPbdepoaxxTnx6w3Fh/Q8xnX
AYhXd3LeN84D4WxfgBaBZs11+nHfXfOIel+f7pmp4Ya+HfC38QDXbnGZx1eYvnNxKEIKBv6CwvzS
mmDAWkdGRB1NoHDrV+jHgUEXsPfKYfsSm6hXXTSVZEiPduFDKOXVp3BQFEDkydQnDaRY3wMfggnJ
OEiPPhsegZeEV76GkEUGEirIHpGBJpBZTQIabwx+picTUbnxY6/11uRjOfmqNRWrSXsvIh3DCb/9
dTRld8zeuTK4Aj+vylRNaAEEw7W+tu8DiQTqAty3Ql+Y/I2YsCJXZss52iHnjl3nVMmNfrm5g1OF
052urmp2pmNegDiDBIDSwl8JbOjHWCL8x1YqsJYcdoMzPMe8ikhK9IR1tW1Nl/U8Tf1thOlRs+HX
nZ1HkPLtFZGFLdIyth/8Ac7ENTcRNthmoq4G4Wnq7t5jLdb0KDiBjfwc8vqxWP18Kqz0g9Jmgdqp
TIx739qHY+M7kqGOC516uvOUL9TMjRhkTvGjK5ICgRE+uaw5EZT06jstvICBy1EhWm9hoUfzPkht
Nf7F5H5+2eY49RYppb9z2nncNr0jA63AoLaebzn4lRH4gy7kJWMbgQ5emIi7ReVbHhsPyc+oElfE
TM5AdL4Rb0BCQTH/KRMNl2ipJHrGV/QDW064qqCFmIJUEetOKvDTlUdplk2tsdftcait2owTsDNx
ivhQvMT1gXSh5OBFealKtncN//zFoc8XANLgcro5uxGfvUuizA3Lup+uHiK+aYja1aiVFve86DF5
Y4vPQfI9D38vBgV++laCvhqe3aZvJL95emts82R7PBSxUzjSiZam1WFAs4dKjzjfDtiWFAOkp/c4
FZ96av3oFPHibR428VI5u4m1RR8DTeU2xsCYXPenFZuh5uTq03GXNg/2Q/MWzzlM03OXZNv6ck5P
JHHA62P/5v69IVk1CTL3WtI9fLB2PfvTabgv1hjUiWnS0a6q2PdWkrSJeB2S7Q5oxNtwdzqecast
AiuZvBiMPWFRFWlHF0wGYorPrcceTv1m0WX0zJVUe2w94BmuVr/TZWTweE8s5ZbfbnSmn6cTOriU
RvpzKmb45u8XhSIBwk0REfthwuLZvnaMl046TF5k9CO73SLHoZphLIsCtrEe3Uv592SsdaVtlUiT
4IjoLIDcAvC18WXh2d5ewm9FkXWwSztSZHEiqsaIURE9o0GgwxzoJ95oWG4PzIUQU7yyHatB19DG
BbLyJzSgsgzgWCLbad1Am/EouMSuX2EBtEOow+MxlT4CnkHAwIab8sqw0Fot3FnWisOpnOaYKChP
mt9nDAzyy4NYUmBJLdYOY7qI77Lx1IqvegmJWnC8T8AkO8D2iTCSgDTr2vvQ31pmuraOcKE3fbQE
wgVvZpIqA3MjYw9n9rYH6//vwW7HS8p3rl/GvZBxutNhbaa94qqSnM7aofCnmQTM5jVbAoOOjHf+
ur91VydjztrXmBN2vtLeDzO5l8mItd1s+fqJBbEJZLruFSMejbVNeY/1zFHDW85q+FV2v70CNWGn
CCOc6BcGuUz+f5VT8o1/KOai8+Vl49TG4rft5ZWZkC1PGSkjezOpgLGf2Em/h0YH13jePGMKkB38
PMvWS6NXb+BC0WV9d/z5sbbOcMOX+zGp75KyU3nwwZOBGVikDChEE51xfTiR4RkmzUE1bZj5TyW3
0I5pWMRxFdIf/STf+OXl+UVEb7rddychtENVZ8fTp4m2teKDdJrglOGFZNuePia/3umAcuxAP3ih
9SLCAS2SsmUdJd9pmSqBX9IYciOENxl0ieyPD22Z1DA2Y2lj3wkWzIasl70nGaDtZ+Uu0PHhoEmT
yHwpMEw8PIoFH0lPdJoHQcOR0MQYnpsdEn3ModxL5Tbu81PWcWZgiFDg1XERaGs7Ctg1qcL3YdpQ
PAjTIbePNJybhdMyndA48zq4aG1SPaC/mMAGGayyBSvXl1ZSsza0ezMJaJQy1xoE81OmCDjxc1um
+wSoqqzTjqRE5DnjQ7DOT0O3XdR4Y3A2jDc14ef0zO3/O1C22/l9MxZ8T2iwWUwU+Nil/dqCmbSt
IOkItr+8D4XdEE+MLuU9yi7L6Ve8Pxh34nRIBhnO5q9ZsLEvWsZb9NsxwdayhTx0LxhOaK/eVG3w
bNgtYvr0XN5yJGr1ehHESzSyV2dZWQC+m6oKtEnrN7cYBwjfdVBZSlKHM9NPm5MYs1N6+XY500kJ
BzwcyKp4almUNCt0hjLjtdXiVXj57qzIh+Kf4W0Nm3ZVQBbLMbrn/wBpm7MHtSlneay/smUHJw/G
b9ZkDCYWok2RC+MxYs4OxtcF9PNF5U7pDYVrZOouEyosN/zeFWIu0DBvR2DiwW9Mx4/ZA3ucBr1h
9mvmYnw4QjWHRjtNwleFvNQ+CEUjN738bCjx5q6/sGIXfU5gpT8VjoL4K70B14OACjWRJsBcBD+8
w0zMTAbz0Z7HZM7ALmDglDR/judKgQbW1uxelUMkGgdMsJpL1lSb/sXjHEQMX9A+l0lB/ji+7s6z
d01M91ZltESKmg3Q7q2TGSu62PBr5eoZqdX/K/+QoU+AReVq2tsrkmW5ojzYSs1m3HfG2DmvB3kG
aeDwRCb7wH6FrAazvcEk/+ImuobXkxvM8IjUgO8jU2niJz+tpvsMTczUNyoQKEG8NtUJAGWl9nfX
CYPnODKUeygnBxr2tyMJyqoU5UCY2EA7Gcfrxru2TJtHPrCcDua51x1d9XCsCcozm733xQrmaCBE
mFUyj8xp/yv0++sABX4QgbnGiiRIV1TyQjduHKdSZhOYuDZxotY6J8EkB39+aeW9/Jo1Te1dKCo8
2wkoHUkvWIIyR+VZGu/23lii5i3JbsnhBOgKd1LMi7aCtAIympIMDfkWbaV4eihUalq7VlfgpKQ+
r+6a1YrPIoBB93jgxtk7Tiy6r8wcrKSYEcOSfofp2s0Y6QkNSxQrxGllX7CiNvms9USCbAg4lvV1
IR+CRJyIi40DzFCge/brJPIAZ0sjJcAAA6/qaMXMr8S4ueiklVKY73iafOtemtbqT2tzPvI7MA+l
G1ubJ8GWBTPzr4TGa7X1SbXUYoC6fmsyCq6HYemtzj8RF/7jsYuI/H+qWJlC7/fYFYbUXJrwOGvb
zs1Dpv+FMD44VSWRa2AcKe0zydHoixylBiaeTCulH9fdl3xTQWuJYuiQOV8R5U1WfSbVxPAOandx
1ZEXW1I3014ek9hqWZkXG0nOyrstZuFtoEC6+UcqzA7VkHxhDuVt5qnG8Fg0SPlGQLOIUwP26EU+
at8O0pFUBQ1sT46gZTq89jybcCYnkwGDCBi7uw8MBQ4aNqw+5ZRRdw1mOTg53BeIkE+2ndbP/rqw
42ZpUgDHE7LG2PjtnZIqFtC9Kj4qFnNHS6KQxQNhZP1IaaDr91+1uG9++1R613RN6BlQXjKJHNjz
u5yJ3GZtQwpUqn/zWEEXgDUKhgke8z7NDs/wo1JCt9jIEeWeYSAp9Rmh8kwhcEAnRD5Qk0DA6IMH
XIdOQ9RMT+8D4+psUffO8RlkXO3lCNiciBni/sTT4Rt7sDCANK9vvzdbDCQzC6oyvHZv0NdOyvGS
TNLNvpHWNdPquivP4lPuicNRrUKSmWQLyL452quoF1PKcB++2D4wVL2+Yt3z8MJbEOQDrRJ9PrWX
8QzGXjsVWw1S20nsKJOaApg1lZbQn5qz/xUGf8Ih4sl6rhUosMw9KYLjEMIDQda3jicHxzVQwCgR
m1je85LZKi8M+hkzKHAbSJiZMNCx4vMBMphy1CZAnXoJuWICobp94+IbNy+y/ExgjllQMRhdw5yt
L2Lg1JBQ5BQBogICLIcJWtjCD40DdI8O5zhj+K4CVeUag7aDQM9Vwbnn3ZlrprncK+Fzfy9q0hwn
VMeIqlzUhjcuB7k6PnfNPNXhO5t/6w3tL4ot9BX3CyRtmHLC/lDMxG1TXs3mcMGxikbpI6dauhXu
bm54mWUrNk9t2OtqlRXrjMGeCHAepewduVkRqUI8F8oNDlz474m8hP0GURjadlBTLCyiUloH+aZA
AuslhQME219N8/n+go+uS3qS8yaRcaf4cTG9K7QMar/pAfWM5LN6+qeLdPg7L1YrQn92seVhtDDl
YoIUgTuKOYE/ZU3LpjSkbK8Z8dB1LGHbl2RdHosJChBJ4/Yq6vwpwjlvzEYDAdRcfrVC8OkMTShp
ljAd3b823c95vKeOswy78gK+ogvnFsoWo0k/uvn8sibfKaVX969orUt4G4SP6UMU1PLzT9wRUM89
ZldGh2wIN7Y40hQ7r047KXowXFX1ptzUrp5BjoYArSIpmqy6dhP2Kc+3I7KYco9fP/LQaqWNHURp
7zka7Zeb/EV80YU5zetBwbOkLkqs4/VTJJsYhtrP9oiU/5O0xoibyZDHuWbh91M+/eA9vkrvBXJ2
F8Cq/4LYgdrlIzDUWr/ZBu8MZLAs8aqqJGB5K7OdC5Fj3+T3wymmHSVjNA8D+TxviXn1ZbXIxekV
/GbSeU7mzGu/JJPT16oPt+9HgenhtOSMrcleaaNhOeOHvScCyCf9AL0eRWjWv2mdIGtp5dcL1Vw5
UcYG6HR1aGLpuDaxlMC6pKS8f0+RkAbW3LXxJCZ8ONcD1fKU/S7f6XlW2OcACsorqZvXMT7vAzWx
ixzdnM6YEN/9DIJDPn02nY1yfP6DIlhYDpKWhV71DQGyovQcr6ElCLQw5bFWTq3JFiy1vIZtshKu
jb+gxOqqaW3GrXmML7TrXJXF8Hmhh9h004Ekvbj6ib3QGG2oucW+4xfV8eY7VT/kUEIDVYGBLn3Q
Uy6rTWuhJuhtIQGznFDzOCVzymZKvWIHVKFDoDdTGArWPpzmLBaOOOW+xVoPbh61BiMYnCxsMBW2
gbeorRAlfXfx7luzXO9SGA6opuN3+BYtS4jBSB3BNOoNF/UPnHYGG8hL24eqWairXLbnJqWkcyOr
s/F+3IhTJVtGvkM7kpiSgddfy2WmgSzBr9yBJPODN0Y/P78kWYegzoVrYS8s7xJECni0t0OcaORQ
Ou412I3gVig9YpahrLSXR91RgKUob62q6dB7fTRJKC2AJB7HcsgiHghvdqg/DkbGducYak+lGJXQ
BPuq6VCUQn3kDipAhTr19+aGYfbxHOWQJRvN/kwuSpxSLLC2xpxXnzFNvo40xecbaszvoWKGTCwz
0tF1qzk5kDxfpsXm+QbLjacSKV70x+kxON/dHioE24FAmjYRFnX5YOQG/Ruo9qMPuA7+nZzof19i
KtVBocKI7pVEI8stoKxUlEdTp6tOMK58YJhbo1NO6YFGCuMy8pkAVoVece5tTB3kkKAcnwWnoU5/
9R4f8JBNdL0yKmQSb1KlCLbo3Hr0zrX0OFuWM+RnuZ63p48AvsoQ4GGnl0Sqnh3EJrMCabjgDBDg
t0OeSQ1mL997VKm+YRZOvuuZdD08vUExBxUGOS/z6uf1EYkwnUcIp/eZOKEC2Op3sXmYayRCzV5S
m0GqOcxlq42/QhnQCjZhqkBEcnnr5Zrw837KQvSv+oajV3Gm4zaJrqJ8rFOsC9dGb9vj4Jooseq7
YuOdBgwPrWrxrctMA66p+l3S123rwZWCEg2NBZoA1twsKv2dri1jjm8Ghyskno81J9/Eo3INGqLh
Y/As9vc4qER3mgJbZuOEX2mmKYA29jOLriQDeBqXgxmhcxpbsNEMe5JWY6chSTCw+KCRAkRTkD9I
EkC94a/ijH1vV5tinLH3N4urIJeZeRPVf2QIWOLFSBxcVaoxdWfE0gxT0h3zBRUW1sv6otgWJDnk
u1vif8Bx3qrfyaYPkYHqMQaZyZQMb3zFUOsfuNisOqN8Ty/ajOENMry7eDHZcw3nNCcCgvrdgk7S
HEqgzrSXnrGWRpIU+X7Fa2+oUCj20XY1PxP21BMLLEJgdO68HmJmPs+GstDnIJ283fN9W17h0eJA
6EgsISg/VoMwJQtI/IYsJUTrBqdDRPATioTfmpQJqp1UyJRBJIqngQy6bbPTJWDsAVMPHRARwGVi
SVDUKHQzmO1KOg3oiozmsqXdSGzJnaPg+eHy1s2bs0Z2zwUYRRQhpvVFfZLAyynxQ2qtbsCE3zEE
iQEMr5J73nh7GOpKv6tEOQUQIM92qLoyHXIAtz0kCvN171+SnOnnWG3UWeKY34P8YKDy84R3AcNM
1MorBKNtZdEHoxuo7wVLhz2Z6VG8lGjp9MTvBPs1Np870Gu8tHcG4F5joIhh/Hc5NWcn4RPHVGoW
SbuDk2w9v5iwl1qSMDjdnwb6mo9YtNiugIW5Py5pPtpn19R35uxMqrVsYDMZLvc6zFX63jS1s+lW
qQf+Aiwajyf4TtTjSUettTW567bgAipiKbJV2PDMYWs9/fo9YaAFwQeYED8Y0HAr4BBohZxxoCQD
50oItdeu38tWRUtuqVvUglZPVU8Ql1gXqSt2AX3bJ/m5FFVbAaMxAUUzMsfEZppx49bncyhlLZrg
6F8s9DQ7V4hAhbAnFhDaSRn7ERr45nbjJ8lo+SgVNAuzJvQ5AJKA3JmDlT15p95X083TNgYtQwSe
jEF8V486jysCpekV19HRfRzBegBCzMiwb2cRSJ7RrAETXhiRxM5k00RJ6ujFheCfiFKNaqMWYPSq
VQBmg6N/zJHJsbGXXLXEc63Trp3+u2XMNNkaFFAVajMI0057ddBPZ4+aYfo3wB3SQ5l22mcZDlkS
jlF0g8v41a7sYyH6U6akAaZCaAuT+KOq/8ZNAcvyI3fd7P7lIJNDNSvi/exOgaiwaFwFnP1CQWk8
cz9HnMIcAeycAkbVXt6sKtxhTwlwJ1ycL5lcOuQCGdOc8PIFYpZ8T+OMg1+dbnkHyGISsVB0aq6I
TtLl1fJ29b/FuNrX3svVVu50SlK6UKGoLMsCsObnayrNVqnBPyHU/C/wEN8ZvvxAG2BxhsUQu3+N
WWFela96KcTSMl2hdAjcgaRosvY1Q3/Ccen+OyKHRMSH2lyxAzPI6Io/1gA/C/JNInzs2C8pvLva
OTGNxT9y/Nkdl1NbQ6X7DfWQonpDjHyZcEDKxGTsTFimb9vopOUdfPBcxX3BihFdBAwagZXV4Q/0
L9A5O98wzYvcKyVEoFdLywlWEDdeuOmZSsntqs+OaQU7RkoWtQMExFK4bDjj9WPqcKfEwqn/IPOI
Vs1Y8xCT3WUoeiEi3ULfisr0lKtH+2nFUsEROY4iCP9JXZC7MIMDGX7hmZVmvDd5MMbqnDsYcJW6
yTgP5ZC88p4fjOmhgzwLCv56hf3uABj6G45BoNfT+qYUedsWxiE+4CAlaiZHq0dxrCI1J83QpR2l
DCEh94IEoMm1kT0NY5z/koYN6VIOrqV/gd2tACu47TYhMAMZOAwm+EQTVhWWCH4AD/U2P3lFQia4
Zh7slD/zUH9NJamGs/RpfZPGu/862al+W0cGFhjK/QXS35aS4mbkiMkmjFAQUoKIow40lHy9gL/r
2QFvko8yn6T0FloBuEoYUKa25mHMnXrefQ1PvY8BaU3TqW7sKCOGiCDRAZFVd8quWO8xuXDpcx7p
3Ipgazmg1Q1DUENgGDtf5WYU6y18ftz4cC/EwPUcDBYCD2QkmwDxWm5lHUMEfiAWUEmImDh77a3i
via4jZumhrKfw8mwCHAH0foGnVoywo+h4TkpYisxC6HHSIjN9MncKNvmH0k2PL/4r/tPadPxAfEM
5TMfOPYR55dVykAg8e2/ol1S1u/RhUnZELUf1ZSY6KGyasta8Cf83i7zP1vZHp4IxUMw/NxR0Exu
8x//yjEVySmKZkG6556+rhWQ5XtPsQYFEYXOKDnJFFB2N2iEgXGioDz6UEudP+Hqmrjr5n5ECxNL
ixid43gNHZGQtyRx0iqLpw2QhmtIKOP+gFBCNLIiZtlpkXfZA4Akx5Zr6g7qeytSsQ/u4agJiU2N
SmarU6dxxIHOG7twSaUfMGz3l9z/Q6v5LttO0cq6yXKqJVVCyUtBAuKyDZqUfaYGORf2/7IdmUn1
kDku+ylac2rdN/voOYJGa/C8LHPFZj0Row4L3viyEySMm8oCvg+EOIMitRyNa4NL7EoqqdGq1IG/
XV4HEPgoylRL1oyl8c4vLIUZhfBbwL1b4X2K2+2ppjZj4lmomH2Us92lGAqcrTZZDdu34xJ8j0vV
ljRzbhPL8hFXAaKs5jHaTvT56p3I8KQzdM6JSjDsk1mNs9GZSobPk4hU2ZX84huTcwmYiC7Ukdiq
1KZ+cBshl9svjYqgLvnJbbpuD4apAdssEn0FKXN8cpbjBC5R4eQfvlk+XtmWfT6TUQX4eyg/3cjo
XgKbK5r7Wim5ApdMGnEiXqn4xW2LntKZ6na76RWxbiF2zMoEyOEFwwVs5VoHgKb/G+paZM6FmXG6
u49nA4YltWeOc5knlxQ+Ac8eZns4usPWAee48AkKeYxpHPJFp7BcLU3eQ/e+/+aAlk69OnJHbQsY
UehinVIatS+YVRZTbOIJ/bch70OdRG3DQQ6PfMEOAeCm+igjpNfw+MFH2ijJD9YCQEnR8FFQMrWm
Q085LZ5WUvL1fCKfN4PnrQShi53CcIbJwNHd8L2+LKyG4+q0YfTMKTtA12PUYw7+0zO1tpAJ/hnN
4PwtxxVc/+7LbUjr6jWnwmTl0RLrlDPg84okixOcmtFLfdxn2ixY81yt2vVuR3U//3vbShuGP3xC
acYOVUXjcgzzrTEX6/x/DsIRk8pfJyuojkBPqTVbsTVWZrAHd2bkpoGX5HdKyODLSGVo5R9KGa+m
RoYxRB5XV2i2mQbhg1ZY4YNufy8vooSuoopu2z+VsmIJkpeu8C9EzE9tBV7eaoVZMhCWYzvJLj3k
wJKl/5TvXAE0FEGobd9InfRLvQ8eR/yraPJGaNIQKGQUSYrBSoRR8fj8Vq0OfOeWtGd8cQMT6MY2
O8Pj6NAYK2TxYIA586DMMOgfkLbd4ZyrqSHu6UsgceJuevydJGhHVj4o+cTGwNnli4T76LoCmEyP
NIEGYbRzQGgmpnSQ/iXoaJf2mK51f6WYLd2rXAP6AnRxncz7blCtPD9ERxtzBE4kmOpW8v3cjd+u
CInrF8Cmpn0VbSIfirYfwQ/KwkSAW+3zovtxyxu3APg5kWJkJVAXZ3ajEpKVSLAiMbTTjvNw+oTA
qYjxBT7v+NhRZ5805OqagExw8XYulWcifbuCKFEmBLM3b9P1u6vltiUyCXRD8FP5UXfRuow9CJH/
0pPR8a3nNaAlJiTzWoBuIUH1zz7LolWccmKB/vrevt6YWNk0YIu07DsjUboRlUKogOBVp8On7TMx
G4uAFA+sSNbU10zCGvHavZHk6NQaZMqRITmG+qZW5d3+t3FE8yPtfvAP25OJ0ckmqTEcUWEASxzu
XtsArsnU/yqg5Rrh04Vv+TDKVQo3qHZtRpA4QYvG22a4oHk0tkx2INijIsayS2YbVgpnLKm5XC6e
Kmy8H3GWDex/9PUJFZxBIcctcz8gIrwjjeeF7YzsFybc806Q9LkQvz1IUvaW7ncE58aqP1jas1AV
xZZ54Cnu/nB7dGjHcW+3Lu0m2mFcJJD3oux4T2KK2fnv6ICKgeOVRuOfvBx4GXhiOusI30INR05k
GL/hTi0nLytFxKvpkWHyWxYdfu1yk9ItaAhnyJ2Yq4GEpPozSHUkToJifNrJmyIyNWfTEINqIOUS
RBlTOLZ74Iu6fNv6EO5eIqMppZRWutdhkMDuwaxRMTK8h3YFCY8/MwQ90Qs6K8sDO1GYYeBscK2U
84+Wrsg/S7QE5p79GvdMwREbwVNYnHmDgBVKEHRuVwltTGJd1uF1uPYprd1zFOI0hocqAimGI339
UiY64nrFAxqSbjfyF+wPpcTb0n2yeZ+RU/2lXDgC2/wylY7/6V3QRcEyF9wKfnNYJOJ2JQ6xFdIN
vvia+wJyB9xIDwtzDyRhDb39dJqT1lbgmDXU85mBN6h/9j5xcGPW4yAsY5/2DHl9AITtU3DHd3PZ
H1NbKrZlS4Qrk5NT3c+Z+yGSU2DAtEHK2NbMOVkZjEs07rSWCTlKZxYEwtXNOWJatHIA5TTtfVql
iqVJh5x2G7taGt6KorfalA74ylLqbn69ZqadnDZv1VqD1UYR3R7N+1HFaVu7Gr1N9y34XBPPj8GJ
cjpquu2fJZpjCpPIQO3yYXT6vJBRwdy+ugVIla7bnn7eM4D9xEI1Dix7NT2GtTVy4keNNnp31X4n
SFtS77qK/Z33r8LWxj/CHaX88fsYHGix/JMpCuxpSwdOYnYjynOXqhKcX/zdNx7b2kaOS99c0mNh
1ckfVDnAx0kc2F9AxMXcTMte/Tl2mNEyutpFYN8HGZ8HqdvBDBGxLjj2gG9tuZTld2oJOLgpuV6z
LZQJ59NJd0PiwrRfXu5qiUzTbyOEn2ptPjZIldLZ9t1KZEkBTA5nDG/sAlw2tF8HiALxQDh5Gmj6
nifpihAr9DoFYdhwe1S/4nPA4zXCgI7UbaGdOp/7gCvrlKF6FmLBFHAKVPxfCujYpQleA0sgan7G
FWEDgBxWDGk/1usP8iqC+HHteeC0K/Lj2Xe14OSFdGtbl8pKRfFS6YjyyqCOLivdLrnmlqR/Wfjw
EMc2Z36N+gBgMpsnZ/1QMoauWIfLAcQdfsE8q6ikombG9JGEC3TYBBJiCPirxeFMfz5rhpo5zfxn
jKhcyD+eKUcmJOp3tXlt37mpkA+YhjUWCC2GYuoT9Kn1sFfgI4YfBhnYtz11bYznD+AjEn9qY3+a
qAc+qG24LOccqvd+GRP3QyY0THXgaIsNdIltDO01f9vrsZ5/1wOpe79v9v7QSK37gmdDGAeM1BZJ
veOJWxYdgu1jLZUfh7StK3O88Km54ztKuRcuEbnYB+0ruxK5VRodAA5ufYHYH/yHHjYLl4/ey90O
6tqM2s7O/wYIKd9dNwqxxl9HlGOCocOPFsZDFoXQ8CqYecEIYX887o77yswNbZDeRFf8tkiraD2a
1acyNdPimrFM2ms+Rkef6FeW5IErdEZWPATstPj1CbzrHK2yllEwUDe11nS3+kWi8jd5uBDlmo+d
zn+QqN0Cj2VPGPKmiF32TB1AXQVhEl/xYEl57N7qjgoD9dRFqEe2q0Cq+DcmfPe+LagpTj7MnAFi
JpK4PGWhTC3+RDdHxgvx2Uld0dQ9jGQi7rYz0JtfVNLgb2LF0u79FujR3AbsserOcbKja+qd4qaU
BZ4PiDntkbqsj7VrSxClzV76tU01k6I8rNyS9nla9gjNm/hiEG6Qys9qEVg7orXKeDSsVBUpmuYd
SVxfMbunbfKUbXuy6ODnUymAbVposw4+9S87soQMP4cJgWg/BmWYjMm5NYusVXSYIn5qiq4teGf9
AHn93qcMCxohtC7SZiQW2uHGAF0pVMUj6DdQGv0/PyJgWvhHP6gVR2TfJSAFwGUqTlT7d8/DVhng
5g4iKQBnYQc0g6eM9Rt2rckUXdD6j214NFmbnXVm5lWuwq7TZnqOGE8Xy7ygxyRalkbYcDe7hPb5
Bhj63kVhioeNMiGGJY9wVmzCvhZELmPErExKUqrawl/lEgMsaUM2rDIsDyYmY7oXedE7oMA9AYOV
jBOysTgHgFFu3/hJKmykTBCidlEk+4/by2X5w8VLlzBG99PTe221Hv/rdHbgLf5s/9LcV/0be2JX
ho/d1PdYH/IOmggqySXNqWCJVlQg8Asx3u+CeeUZY3FttR3cHHcZlLgkf/qzCDfrx3SMvMzSRCuA
k8/Pb7QvvVBk8CSG2JQuFTPaRTh5zCQeKdBbRRxm35a7YyfsT2edYudzqb4UrKUQRG0XfyLLul0n
019SGyO2Kz8XkOBvzkBV3FBOStszWkkwCA3HjQKFaa816bTd1ZKL4kB4W6nPSkOFcaoj/8Ihvo7J
ac9Nsng0sX96pm9opjAi7nTkOFH1FmT49IOi3E72oijFckRpc+cfXL9RF7ch/R5UHY0UDJFEdBEH
+yT5C2XOrf2V+tDxfEONJZvVvGBxqNEBWhYFcPhVuEqQjXQNqBEhojI/O/9oZezY8ldpoNQX4P1K
mPx6rx962vxhtfru7SCqrTC0k6oaQf8MCurDkDxqU8WONoWEGyuI3xwLbRFLoxc1JeFv6oiAkxEr
lh4nHAGWtSynNqkDcg3ZNJ4xBnHbh4E0nFzHrymaY1GrkP5DHic0j0vlGfKSiAOJBmDxDHMZujEB
aL0JQNgfaTCi8eNfL9mglWcnoDjLOcy0C7+OazaBv0sNFmsNzK4VdLAdMTvE5Q5Q8rneuSqA9VZb
2tEbF02CeiEDc8vrSxhmJ+dm3K6yUvdR2XGWDDVHVuk9ggYcu7mKXFn77E2eR4TR8FTSk1dUXblq
QnvQIldSKOfSj2dmDXpBoqmDVvS2DdjS8T229lZcGhmDHL2HuPpZgmM5j3OATuRM5GWr7G4m2xP8
G7d6FGme8sX1aijkGsobyjPDkiuyQU3ZNyj8NLKybQVOCoTfQy3FHqJ/4NZyCBQN1+JpDtCOYnnK
Chtm3UIVyHnu+OwCyw0uOwvhjdPO0KOTM6cxY9BZbVCDpH7HtOIfxD6JSm/ln2y6jUkg3l4TeJtY
OJ649Oh3CwuCmks4r9W6hvJZVIgVpqkotc2ZKgRjheMCsKrShZtL6TdIgO9yvrAtmU10CKb7f9ui
vMj19upM6LxKohR8wAPiHqO7GoWSJiQsffuFaXpuxz9W5K2PmMhht/271YvY8Euiw9KYk/CwXfcx
W7yyyiPgNJQ5cSP+zAgEmPkt+k3SYPQpsxFIKVrYG196KIYCGM4sQRCS2Lp15TWk+zla/PyrKijG
w+XNhULBOykI6ciemTECj5cCTegWyxcIITTpFpXNww24JvMwyQZYpyFvyTQOF9Hi2NncRl7N1wRm
y2jX/dQFzcdfKu9rdf5tQ9L93fBZSkYLYrblMo3VTPXqC8nNuIunjoSf9pciY0fqWQmahrKLZ06f
9xpHE/PtNsyJJlC/T4ro+n36ates+/E2cG6BAwDuoxlTeK62dPKDgVeH4/TTeDPK0QSa/gvEK5hU
e2RSN2TtqoyCiaautOnzORO/YKXRrBC5dkKzAOHU6GfWZaKiMksYs8e7dbYLAZR5NrhSKwyOe7vc
iLdY7BhBCAmvv5rUOx64ORYiE9NVHt107G0UadMs3Nt3xOKQvWu8y6aKuGc8YpIXlv/yANUlcB7W
6J3C/el8mTMS9Wu336bLd3sqOqL1ikHk8WPtxtvthZfgkvATlJyVo+UOgQoqKAa97c0KDEZaIQxv
VtiTyg63X+pYsyDVo3kfe5ylUhoLUHIHb/jUs7QP/uSm6ZQpCkxEN7XftccpRzV64aJEhh2rMvwY
GfbXVcxvebzopM79i85B4P4U6qK8m2//sSpqNA8BkByNNiYjpV3/PN6Vn1vabXbYp8DbElwCySir
lEScSgt3ajOYdJco87od+n2IxWOVaRionyPKywtOlGo6HtVn0zl2y9afP3RXXCOdOoRitL7Wv9a/
dCxdmQs/6k1es/8l/p76py+d/VFzDa3pBk7agxDq1w6sPkRc3/hybJh8QlXA8Pq5cQjXWI7J9XDX
0CvPEAoF+BXst8bSbkBsbklhmXVm1oK9BKItvAZEhuc76dgCXltnRFQIsrH0CewQom0UPTKomlkr
582nWxvxf1X8VfBzl4I4vgK7MLLfMZphCiReObX8sPrJRR975XpQ4heNEc6tIxrXt4EVwaBLKM9m
48RuA/zmOmmJURekF1LjubgGnA7H7dXkchPonIcHhCg5qYa9BD7ABkrq8fOs1/6EfX9LyYKqAM2O
YEQG4GhtzT18/L8LrTRNqjgEiyUcYSVE1hmgSaorCv3/Lz0wWOg8sAAQCm+0qfprLGYLmAJE/v+B
r/fifgsxWuVjj8P1Uv4Yn99KQGts1QM4hiVBl9Dtg08fhbh7zA3RW3rSRqogdbn2j4fpOv2IpgAy
s3dhWNut2gmyRAk/tKq5SrJQu9QTVhahAc4yUD1r0pPUcuWMg8mDOWqCS2aPK5JQfKvMrWceVnpp
m031HWJ2Lr9UEtITqyqHnQuJqrWB0F+uHirTy8HKDhASynLIBKoDe+y3QGn/IVzmERu5HXHAwxKE
sVKIDUeSD7jv6ukvfnYHzeqprSxKs8kPS0RTDQdRew/Q0qtnLPma52O1dtn2A8FyaJdbyGE8QjsI
R9jYaBDqQo4qdd5v4k08XXLVQQ7F7wSYFD6yo7U7pBCjJA/9pfMKpdMBVb4FQdbB4LjF6uBPunwo
NZ47K8/nTChOOPq82VvYvFJUNvOde7KnOXsMlwXcWNTdEgsILHaHmcX9jGScN3o3emUb/QQMNF4m
hHPwYoIkph4byxK0rAoVVSfdwudtt2fbO78OWWTsCBpCOlQZimTZz+JHqly6JxVZkO5/zpul1BKr
cO+2h7dj+STiCWmR4kmN0l6twhe21ad3EZSkzz7nsa7HMM5dbvYmSoy0LCZOBt25jNJ1EKJH0n5R
wSxkLt7iSXlR9sTCXQeuc322mj1rkQp+UwXxA8ayy2b7zdQcvr78Rs2Ugr7ireZrS0E7igobdA8J
bi7x3Tdj8QCPt7vZpVOUsVApQxfjEGmLs2wtUh6PKkGWXzcLbPDc1XV1+mPmFaCr9aNSxjNPZLrq
KM26b6XnGCYYdwHxyyaIRS4sfZ+k7KXRvFrKq80lIDQfAd2PMGsTZx6WEn+/s07BUPOyjrN3RF0b
M7cKeaxvMHcPaiKNwQ51q3d9FwvYLeyJrAS3URfZvcx9RB9n/sbdYfnLzWIMaI8IQ2N9vSB/finV
7zNTgL1J6KvSImNEQrxQ38NQE/s+YCAt1LZWKzsV63TzYBcUUtvfMjbhR8FKdwKbCPUWSnI4hqsN
8r0liW2H8zbnU/5u44YL+NRC1c2pb++1XK4AK5D1zZ0QjATrwGqSCfeGbE6lzlpEuUCfdci1KbG5
hCRT1qdUcUzKTVmu5RolQJhgvedWvz0rfI4G8QU+VS2Pl++O8EQnCeGGBV4etm6AkoXqyfqT5l8s
aSg3LK56aot0ka8wnDyXiDCZrTSFcIQQzbNZsESrA9lpHAMxYSvEMzACKAAwinTHEGaZeh7GTDKE
J1ulkuDO/c1GHF7Qi1uCiZoJvpZKL6lb7mA9c+sq9aNPuigRFUECsxxFyWnZpFgm8Xi5GpmG2H/9
lwo5j03mMwHWmC1UkNfb8hJU0G4pIpRnW05HzqIfvAIxga+XCx6/dVaFWDVAcJ+d1v7J6he9nCcC
9QSJ3yLTe25ee858Hsx2a1m1tdqUgaZATFCTt3ZURWu/0r9eWYoMzhbCtW2VUqR6NaBL+M1vrqQb
qaDvgs+f1RWpdhCLJld8l7l2DobBWW9ZuLERUbzaBdZJiUvL+atuTQ9o79gNFrGlqNXUD+FiflKw
GGUWOYb0ZLAk55x+1+mhsAKd7BmhNEsL0rmdxJZJ/5U/BfoiTq92A5YY1LJrsP7Ye0HcsNO0W0mS
hyjeRA2CMA/Fm70LNe48kH9vce2ingY6w9JdE01dsCrdzApLg06m0iVCua3lk3L+kii28qScz2XS
uBfXwTjf51yEDNRIBwV58iAiDirT6t55dZ8zaReEZ/6BQUcL71+KYA3jFqy7L92LeAUKpdhJYDLb
CSd+ENBbTMPltlM5nQTwWwJOJYQtupJpeIGMMGruwhvkF8qqRs0YO8pjXkO1cgyeVYqMwGoHiH4X
YnKOs3Jp0cGxf45r/TIr3WZuOABh8oP0CBAEwMG2kuHocyPm094bm7+hGVSf/z6F2vltp90hD0Fx
Luvkt1gWMwD4aS9Z0qHl+Zd6oIdUcrEQ9hBrO+ZJ+qeabIhvVaN3xC2Od4zK4FYRM2eCVW2zwzh8
eK8ODsSS3kAzQKJWEuhdBEYueWupxmlLre8mIGIYpUtAhMkvHXGTTMBdHJatwVbErFUSLUC268KQ
IMdU+F1xBMoLltJKjA18wA3uTaXDEU769jwBI9ml8A/52i0/2Ue4sMHKrKP56j+uykLZSOlcwR+S
cjHi6PO/PLvjhnLQMg6dvhNQ/mi3X20ZNdu0wpHHGBH86DovsE/cfVF+UCuE52ETVSMH8MQZOINh
K14ZykGL6pB2NrfQcBJnuB+3megk0RS5fS7Kl6JS8suP/Z7tp0O8sMdCpt5pVsJ6T8zgXPq6K+gw
3q6KhDyDNUITIDp6WLQvnkpj0pR5Q9l4w486+yOGw1cMqDKwMF+ZNnsOsCZ55oYIqe/hJ1fG4ve0
grXjVk754G+vHYJTRDutgKPEUiFTF/1xDkvMnqOL3gi8EKEcfUdyqndBIPcqIV3iyjbWXPCa/F4P
9Yo8iP2N9ueaX4Gz9bXUtzO0hynImtlpDzQIZe9bNsPtwCObeDsbMHMagsfsZ4tG0+bkBRxhJSrV
ajUrAax6rs//wasvSNf0WDmWxtJqWpZGVR0IwXjykBdpC5wq3Q4C1C1luZLCCfmcABt880G09aXR
nTEqCCm3Y9wX0r/vI2Rb6b2YS766bpmh8Zhp+mUNfJX+QGYOzezWtuIhyQxSL4Niu56xseug65Mn
tZw3pv9pPkeQdnZMacuUQIRJbxitvsVqY0QSjIxYN5mI36SwrG2fZm43xisStSfWwx+5FzQRayxf
qV+M1p/BpTPTFy7K3E08qz1J2nRuJvvwiBUo/sG8DOIwAkF5K54RtbmNy/Xi6oMK52hEGelq0rhN
YnT7pXfH/umPPJn2DbVhGyR3EpDhvKuIPjx2ghc2AVCZwrBT70mM5a8oHT2XwW/FWuqF8JnQEpY0
sgkIE371OmMgceuASsHK/UYSJG27AmVU70FWjKGk3gX4qaYtz5gcGLwswC+eQAEH7ACs54YgA9f8
d88Q4nzyZl3W7q9RTkX4WBHTLLOr535wulya2Am00lK1YPu0xg+x+MPdT3aMed3cSUId1X4U9GYI
brvnAPa4UbDtAsbE+pxbO8B60gJHLzmowYiNzxWK7/mVbkJHak/8nTb3lxhHmMtARwWo5cOTgkEV
IQR0vLnHPl21/+EacIWK87LiWk/uKvVAMSX1UfN9hHLvaZ0N2Awbc+fDFdagh7YJRqjligUlpdB6
ByPpHGYIPGYaadc8dDdRJpRzQ/otvo+DUTwGBZXNpy2DMs1gxNc+SypMYyBJbnhZvbWyWoJA2xwl
E0WJe8j2yk8sMgPtnIsgibv82FRkNMWYbpVj2DOc4w0u8e9KpmpZaXDegOUfsh36JQnkYUvACUQl
2bLO88FOmugcJzamgX0MZTbGZq4Qoh1uWuYpzuDewMJ6fhlf3HNrzMmeZptP9vL7XkyveESOZ+m3
XWoq+k1uSxvZuvjlxyMgJeHBfWStfLy4VH1omSeVW/uS+/JUm15cEL/73Do4Cocx/jZNlt3DOjVh
bmmSKe/AE0kzzvuxKWNkjUeAC8Gly+qnLjAFq0qZQqav9Hfsa9Ko1mnXKZ0KvR2UbJ7D0cGL9QXx
OyjWoEndE1ymvCtfJ66OPJxVzUs+QgrGawjUBizQwlMtDM7QSfbL3iu8bCv5+KkIfYHRaGebPchJ
ORmSEeHqzX7XXa8qfdIwaJZebf/SnoKBWACAz6vK5eVlx5LcX4WqIDtZ4X9KwmxDFTHr5L5Yac1F
hDlCDzrOixHC3NZyohyrcOZAt3Eq55nB9+FW6oZx4SPVCfNWzZ1gPiBqpfaSU1ux7SFHt3qRaeH3
EERK3DcAlr9nTxs9nNmbu0oh2FgHyy89FELjL35YlkeoeRhrb0I1k8v7Z6/OUvMYj8VGB+TXLeM/
8+80oclSmIWQNdJ0kr5qVykXoCq35MDO2SoVOhdV7I+MFnfWNkwruj0FX1OcLKc0DfLkL/vAFtNn
N1DWZH6PmYQDXjqxmbjHjqs4hPv+rJoFFj53XFa7BnJVfaGppXTjfZszDbSRqL4/WSjAmfJ9QCeR
esGQ48yWJjyfhSoWGtKNdgLL2shb/nbrlpe9F4xsrvWT3+zOeM2LR2YzaHIW2FzEMAw+qNXsJn78
9T9LIaP5iW8Z0ZthQsskzKfnmyNplatgWMrtB7A/iREhk8kOcow+iv1P0Nb349b6F0FuGD57OXjB
+8NxKBXdrcDEXy/xjKrCdPUikpFWP9Gfk8LVnL5BUJ5YX0oXaVjSdoehMF+jWjn1tfdZIWRm7wIi
Tg644CzyAtlR4fI1FSJ3xaWFU6W7OCoNZHbKMeFa6rVNfcfirdgYlGumQt0uAWKuY/OIXIeabY3b
6HsrVwNWukq0GfujPt/yJ6/oqpjBAC3XGsq/898SAryeZPB1ZKkzk/i+xtWSfo4Fj3evhNUKL6/g
YY27Ci2tXdHEhyTD2IHjDRXEakH8RjAU9zyx+jFRfHa+/9/8T2RG6UWL7IjH46EQB0y/FiWjRr7P
Jkb91OhzTbpl542Ks9EF7QLqm/uVjpY7O/32miVB1qSX1N7g/7AV5nxMHJEAaophnqucdG6OECpF
9PCAO6j+FfEfObkALz4xDkvkvev+R3zfZpM5rRkjYoGrKsPPSUDQMjrTGCym9f/b+q/P8tzr8Sek
jsVTSXS8uDxsb4mpr/bIKyX1sf23wXHrfXwK1FYuotvPk3IGYMj3u2MaaNDALY6oXaQZA83K67l6
mIlnykT3Wb6iMYuv556sU5liRJSZHrPXNG/5pvbm7nFt0c+am2efF9bZsQIz+/CxFXOlpPdp9vNb
0+lWWWlc72FgSauzduUJq9MPbxoxdVEHLnvoz1bHXoIOLf+eqgAH/n0fUsbPztj6ESwmMc3IuwxT
1LN6SS9EdKewwMSfAv6edHueBlzaM6Du3OGFwzhkoi+H0P07keEUwd8k4l/WTBC1us5NHFpTph9r
FdJZcZrfxi/dAYkd6aHqunQI7keJWTf10SgwzrdW5/MbTR9hNbf2ZYgP0fCVHU6wSwjd/JOb2dME
X43FTafEqPTSW+sUTrLO6bva+v6UPcgydsN70yQPZJDMXXTqVOzhWvexXDTa4dQmwSaqD3SKb6au
JLXz37wVCAKRskLuzEt6xRobs+1ghb8i1SD1ot22rK7loLvGUbXZs4mbZdDFyUBFKUxtOT381QEw
nCWNTgAnlvy50u+uVjOOe3i4Qy5f/HqloAb/08EaoVlZbDjqYeaRgBXRQVUyImycRbwkrBcDFOga
2YoL274RgEw/tL1qz3tcZxILcA7PmYNuAyY6VbpdA+OtUGAKZBVI8zocm7xh0h1uAdsyIBTjVJTg
yHtb4+VK28aTcsel1z0mmZoig15opnB1ViJUALW/X0u36JXEtIehf5eF5kaVTVNGckBXgn3SKAcB
q+KxjhydYDWCLVUQV3zmmYpoYI8LTy56NGa2fHsTN9u6Lw+4ZhzNMv8YKoJLYUIeKVDMBKZtEhQa
4Qpv5u792yQuwoIRttZX5RTHJEGbg7Yncj228ZllqzFATqMnqeMUdLxCoSQOKa+XjFKDltwSayvL
EUmc45MYV2Kd4MyYBhX6zOcKxQUmmv7aFGS2sIHzhPmw9QULhpIMEPWPiFATIlB+96c+BCxBbvog
6Gw+yM0MPf0ZouuVaw+2pC7AP1ZdlfTU309AJuAAfT2cVklUOr5NG9rNg8YSx7VPJRMjGDwZBAqL
WUEuo8r8ZIOjqcJgslQwvB3zf5cRhXl9EikfUjZfEfQUl0c2qeTumTuSdrwj9BNZ+Um77PEsciZd
gtmm9zUGQqZ5ZhRIJYhiT7EQR0aoC4H+fbKevOT0CbVJQQfxr3NJkqWVqBQeN45+2wwG9aRYErFk
31GaAiWB11SMlZx47KWJ343R4aM5RW6/mf7BN8G0YVQWWH1E/Fp9ZPswX5jjPMZTHmN55MR5B9jt
vEsRg6tIOxYHWt69Y5mIUM4UUHcvfLDX2UvmVQHpD44D2ECFiJBHNtZk4kq9iDwPtwl/9fuMeLe6
gDABRMbPq7VZlw9g/6oyz40Lv16OVN43g/XhtLNHdC5nT9t3PaJnD3imkAXKBSw8PWHB8fE++FUK
a4AU/NQmak5KKfzMeiFVicykQgPPKOazqKxTW0DiY6nuSo2Ul8lCO/8Ltt2DI5kcXMqobPU8a4Kj
itPnXXsgrcRX3fbd3R5a7c3t7IyhzxWB21TYMg+mFgY8Lw3VtSsB80Yuwymf16Dht/tbQF8oeUMZ
J5s4o4ELqg+/2ICgTELEfTL8D9+OXaTiKzAGh+G7uNOjJkcHKOgpltRjKbUeaVfySx3Oz9WtFLnS
FVfhMeWnuj5RHm5ZefUrklFCT4SjboEpix+xrQCgd6PnuttdR5VZP3V4pUYSWU6/QMEzsx2+q7KN
Ck2/xWdVH3laYdHxObk7marW4OJbzwL/m+Nd81XSr3cyab/pSlM9uKfXWFEp9Jd/4amjN7eQnJpI
+44d0nScVn/6Sc72Jpk7jLe+2aSDmdyLaedGmt+4ngkpmVOVKFkyHyh7lgOQWfnp7vgwdCvuWvQ9
/8oCCMDHcsQPhcBMOelifLE7/OkEzkLSI9aYI06lBUdYNkEbV111dhdlDNUeVg3lIA+G6wrC0piP
rj8kioCPnAorw46GAUxlagIQWn3A5R5p/q9K4IB9FBQP/j2Y0uAFqKHpR99OYSFYsL68VbCYeCKh
Tger0nIodz711NOBAcB3av7n+W/PYI4dPh2GHPBha1FXRvv3nZEWzr3r4+LXe46bTox4zS7EbT9Z
VvVSz6QNXKMI/IeIBvk8Q5Jy77hSDe/gnxDRCoQ8UfSK7tDvjQYWEihn/Wx0F2GXcxhgVvOgdAwD
097QaHbOJ1Z/MMYPAIL1MH1/oOcFc9JB1h/p8tpc0eZgDUjpRcgFYsvlhl+aGW3aEQvmfFKIcSMW
kWcQfhDCbIGy7gHDzPhwdAyEHn3v5D14lHXjop73EihVuGJHo6sQcZGleOGL6RKKBnHmv6XVDYVy
53EkoyL3yPOb0NqLfEc/4Ag8ZySAoQuwwWny/cjIfRGzCntGIiJd+9QzFP52cgH/tJ6X4/X/+yb1
EakBLF3b127LPrx9m/WE+9wJfqPXiVQMUH2KMbGlr3EBGAsPbCyofIftikw1xyn3VONPZkt4VUY5
hg06NFtQ7zoI+WMvqANhWNn5MpBHoIi6FGHxstxSLfwj7Lobskb5oLmI1gLL6DagHYn5H749AMmB
mBj8hBl8mclXXYPHHPMSIsLF3JFCwU+8ltRnqoATJvFWVenOBs2B8fftDLT8dJ1yewTubs5Cmv74
W3GJLuqiiiYEHJGso0onkVvA560nIhBgS7IHgRjDnlf/O/DFXW7aym9oftYhXO8jFb6/yfeQmwKU
NHNW8EbAEQjZFu+mLWqCNsV06ywl05PCJEAyVJlfGFuo7hWPlAN8XbHEQALICWSLfIfVVPqsEGA8
15K3mAA7E3DP8W8Gg2LzwNvWahXcA+B2lm2uYxk11s/dxM5KJ07PARNXKSyiqFnA7OmYD4GZFf08
BCAexbpGIJ9i6s5rUr3PD/Wlelo1Jd6jPlOdxhDlm2079jdAIddJymx/qGkMqMCU71s91DCIvhyo
yqipz1GHYQ3Tg1IFzEhmAsiFkKBFIRaDQyIuFh9F70U6DKZrrsinW6O7GtYMNFJ4MzSoujH/xJ3O
dcGr5kTs3sCc2WuezDNLxSaB0pEr9UEKvNUJ/ueoZzzcV9sa3cYPxlYbDLztJPWAd3JRv1D1yXZd
YpY7dRQh2lx62/Tmaf1l9b9q1qHCmsS5Dt6owVTGFv1kabmW6emwUOd0bOEXP+ucoayFnQ4IIZnN
WGT4xRH4+mU94VlF04Y/CRNnr1YReMObeJJGpW4PgS2fNIgs2LVnd7m0hUgghEDHmPC2OHS9ZbUi
ZQ/wFeWm7v3VOGXAgK7XOC6XpOAYD8rKzp+2yCBzaIQ5y78FVIH8u/9gIirhzU9GVhDPKmjjbYRc
/6ylAb1dBrUvLoUQvuBPZkALqPP8RUn+o8NcBKExtZ83MV510OZ5MxFF2jPn8AvxGXc9+VWiusvr
80uyLIJ3gvshl36DGkZ4ZXHJP/D/Fj41nhH8xmH6GxbWXOhHoSYiGm21fyfYTQ+sM+R/AyzI0cBl
HY31lbLnbjnkPBUxlORIMsmAzHjWy1audGOl1NoBuBBo5IpNSYL4jOCnC7OXZUokFPOcwg/IdjbD
U7g3NnrIZKCudpFq5urN1ETTQNieTTxG3+I5zqjrEf3G6XTG1PvsuIGEfm4YF4YwAXZrpX9o2e0F
T202s9joTEit/Jj4FT3siYRi4YOmrVLW2J2F+PlPJx4tYCqKZ1+1qqdn9ZxrxcQm6uFrF8hpBs0q
qcvvYxbGtGLHPVVAFT/7zeknkrCOMtnhlcQUFvekRLBcO0l0Ec8GgdoC9o7MEOj7NxClDnNpChJI
4fY/cyZTjDSvHLMBP4YlP37KNfJV6IQMPc8lmwfMrg85gD1vvnPtjJwL3Tv3F86GTxoX9oLNwfUA
DOrCZFdv0Bt2+kDwmm5T4xcj8d7UW34M6g6I6wk4+9gp04XG7DK8Q+NpEhWzYVb3LZXrhBy8Gh9n
0PmPhhXa15nCmBOEk8EuYiNY+bFNg3hsjspg8BGeXznv1lfF2H1uP1OnG3+hF7n8hXOB2Taxv6oF
za8iasjVCDIjxQ51qx4I3l6QVpUF1+J1GpPjd3NHtaJIK6l0y0uDr9aDWGmNgId54/hUeUwHgIfB
nghmD78t6cLdCych03PpRd1uoAgQ5q7Qiw8J1ZufsEAPBqU6kBLvfBb78nm5StvLKb/fkgjfXern
FctHwmMXZNtILpSPK0rdN36vKjCZpiN3jFMqwlc++FCei0l/ohIKerQpv4oiY+J1u7lYTr7puOXd
tjicYiJO+mw4K6FuUA/gxwcIO1YcrPX8i/BS3+I1qW0TNGn0T7ilOuPxaycQKW0Kpk5UMnUemXEV
sFAzUNbmGzhZVvnZwfQ+TnVCr14PGMJiqBe1DpVU1oaolenEQq65W+tghUUimgEZyD+9sHs1KbUy
sP7VK8YAeTGNdEriljCm7pCQvBxY/EBovjudpwptdSiBE9E7TtRSPnEEtdXX08o1qMt+SwnKRUyD
cDRkeuqIx73HbhRQ6SkNj3ZBiHlTWbqNLAm4jZwlwQFQ+E+l7FwyQz9So7VjwtpfFyJ4BIEbkRED
aTUSMR83t3MICdnLh6BTLVspVNO0RwuU+3IJyfFl4vGtKnf40KH4cIK8YjMHhWDL1py+UH1Y0lQr
EMiXo3QoZXEwMBv3rNWW5N9lSjwRrQwld6RDG+7N2w/jrO8l+dkd+mUP4/Zk4eJQKZh38H7EPE+B
WkuerCpoQsp5c7k31q+6TmRD+Xfv7TAM7/RKwtgaywHLJODe2foQyYh4zp19y2fRRiOoCmt8dv8L
/As6kEST5SO+43XKMqTMJmruSr1DOpCNpQ7cxSN5VDO1Lemv1ACBA0lJISHpmn50h6wWQB/HydlO
pMkMSiBF+JbgoXf3pLmeiG5RjN07GLPzB21LTJcJL/+1HzYlQwpFsvJbGxrbp0ItR5fFCd9F1rit
e0bobbsTV7dpyHrqrRMIFID1hxAFbTL1qIjzDmkzzp30dbym4Bqat9y1ZW7qvWAtNbttZ1Fmx2KE
6KNmC96z+t3R5Oj5wx2BquyVi+zp9fTNjoTgaAsUDizH5HGxHf5RkUo7MFh13tzuc3xFrcEMeoC2
aAqb7gFY3FsgY/QF3Szbz9DfJZgUl03O9A2T213GlUyB4pGx7gpEWlXW8IR2iT/G1PkiTgvJ3xV6
hbGMaE67UmpE44O69lpHSChMbwemmXd76uPZZJj1dEPp/wZB9/yfHLlgQb4NkzhDK1S37OKG79/S
8PVFE8+X5DvlfVsW+ovPIKuHN0NZGJBtlB1nzOYmowO9sizilZMvj+YMzrA4za8PkxG8voj3Isi+
BLMrRWbE5dT0/zEzi8QVSaPs5QpDOiOEAHhZYCO9qorj35nqs4mi3mmRjx19rEuFUl0L9QNT0DvQ
fsHJiFkMvSZHUaATf0Ok2sV96Wy7sibQ/VoGbkXQ1pL3WN2s5/ezHAQVk2axWKeZE8PduESYPjii
sDKDjJk5lf356cZVUCULku1cI28RSHZLibuxaUCrXFNu9bgjWHboqW85VVYRMeFXAMx95QHPxq3y
VKkhs8hVKdh1fYkiMV8t35EAS6mb9uQUYbja5Rh3CmRh6TicoSH5UqtqOGvY7EkxwakPhtdHVe7a
9cvsrCXceWh+072I6QnV0T4R9qQdlRGfRypIS2WWFIUA/u6Brj7fCPtW1YTxuc9kr8dcfQ8fIJeq
2YbKxIFWAMI37YuyoFmGL7Vm5N1soY++JIJSD9xU2U0KE6N+kMogDVKTtCfCM2HS7b6hqMqgc30B
J3LCqXnqw67ZSbvSsStW619l8EVi/aAy3MKRwoU0pSJFPAiZ/m6G5114OWHRDvXobztiXkOaqE+d
JiOIpn0yX3vBmT5w8QyFKJ4TaAkZNZnRBs9usSQw1uXRbwF5ncXGbFRbFID0tqvVNizmMwSZOKHi
GWUNljsruNtK+x0l432uEyZhCCz3pR6whFBhfT9+65Rk48Fp9CT0yKSRueSBTg3UUA9N33cv0pBK
MO5t8vh+tCppsRBzML2888/FTMhVgT++XSGg758cN565Uw02FbfR5eEqzccQ1LpbT7Mb02Ab4R6X
gFV+QXpwTvPgXT47VdFNcG2DxXfmlSgD54z6frwzyWJbHJTRxf8fi3TvGP840GoJtEZTbuJLc3sr
wmLhToeTHhd6BsRBM+Sfm3VAZihzZvX9QMycIhoK6usSTMDQagsm4xeXsFBx+ADDZHNmtXOEkVh4
bKHilc/9RDuHJyDhia6y9eIoT8QxcJJSNkRkF/M+Ydax9bMTHJuRbFnn2CPEQ5epctX16RDQL7yb
liaQdZgKt63Khrnsod/DrBzJyvtoDLrv89N4yFbAYeXXmqCSQdxgYUE9tPrzF03GmUR/Zd6PeG6/
gTmq2s4h8THwcJPxeNrNr1WTXgta28AYH0EBAUKD1kb/YmxyaWL2MVjLcXF+LQoDX+NEeNZvtEbx
zqoGoPmwe2jRbqBhUE2zX34T2xkpB+j641AtQGQzpyFDdEkcgqehmMnlhvEYBYIqQt8b6E8mfAx3
4vjkV6lhEvZDL9hYDc/wR2QWpNzilTuA8udugNWC+IDMsDWLcqpNz5NzSWpSubxR4ZQNBqUQuN9X
VMe4lfYJE1JYshxbQITDZgXGCA041uZbpEq7X14ToaEFmP/RCIICbbIfk9+FAGnpv4pEWRcCPqTl
pt78EFgEzB2gCGxoOAd2+JGW3Y65/GVJ0yTl04fIE4hfVDIHlSHjl2Cm766TSFLbLUbPMh8uzTNk
vqgIPVz3JzRc2iAIH9RPcreqt5AOtOac+xt60zdZB406jhFpGdCMwjM2SU5Rz94nwiUATRgeibkW
trOZW4Xj0s+7yKkXc82/nYAVycwLeF8iWBNl1QQrCDs4xOgjonw6GtdyJQd1AaFq4L+AFlRwC5TV
ozz6rKNJo6PK3jkzHcRwr0/eaYGt0rI/VcD+aVg/goq/Kc0L4T/Vz/9osIg/rZ5NG2y6nIpDhNoz
rNXXYROU7KixvMWMYJBwVzWdArWyrSaxGNsFWasFQGYs8jmKFK+2hUkzf6liil2oyFmaLJdA5gxO
nbwiox9/rIb7MZGhzJuQb4+27ptfZUMfotgK4cxIRBK866/b0hgvd2j0mxWvK0uBxfMNhDYLnXsa
msfyfCearFaREjZZLyiy2eCMDljoelGuWY6UwIvf9BJd5U6mi3sllZQv927RMX+dxIVzffFaKBU0
h9VMDexBFgctlsfNYuM/yhPicOuw/uMN75eWZiyb+GCIknKd2bCfrX1FbZx6ct1J5Qe0CBqBpHA6
PC7JLlqtZOkBMlV/fEPMwJ9Ck37jnvc7sDzeCqarjwtcpPc+NhJ5FD/T2nfaQ4sPbKtk5Fpk5xK+
MlGa6hR32D/u/plxdL8dVnpIJ4UQ/OKRvIonGSmZt7LsHQRCvjDQhLfVq6UCNNURZXu8QBO3ypdD
l7trXx4s85tJYvihSsmw87UpxOvkKnk3TsIePEDArDwzzP/J5LRmKXa/O4Bapd0NFvDaqjNmRSLc
pnmtUEMHbBSsR+qCUaXCpLpi9Q7gvt1KXaDBI/V1tj6XuiWkGs/gSXn8CqSwEzUofdjUduESd6JD
CMKAdn4/BmrfH+D1dRCXdFIeJwTjc00uI4yJp4GT1mfNKDGiTTWNGLMVps/Q9cTQCILE8foCNFSC
rDz2wLKdt4WXAuvbpeArKtBw7wj3OGyeOs5YqiTDsGXAcL5Szn+71DkUzbjpumbG8aOlPFfe1WHj
UouzZSs0S4cNJ6CHOGhy1YmG602mNfxDxC55giag8tTiLTD4qDeNqYhwpseknt6tvrzhVvflL6qo
ufHFhPXrt3tRW1pDcOAHQ+sZ+4wUW72xmVYNa+TnxZE/c2YR0OF72ANaIT8VHFhAs9O0w5iUmVVH
/FUSFFqOIVBJRPdVNURU1hWZBB9oSUKOpSsUO8rnkMYqGSPUqfMqV3rkpcoPfahNsZIMyzqtqw2B
54QyU7lwqf7lnA3gQ2EQRVY9Jl+RAqZmtVh2XkYiijeP+moiytOiUH7BMVPjCrJkUcjqxQWyHM6j
pylJPZqQ7e5FRWfaYZny+JjGLQgLOZW0HODmSOSg3DUnNrEdiEAyDuAQKqeQL511k5uUt32B4uWc
Ya2CsZOVwGEpNGJFGOL1YAd4U+fSr8DOd7WndKq77Y7bVGABdvGAc7r9aSPb7xz90Dgr4HVP+ZH2
OQDmBjWWyrU4uhhFSTOmr4TJmFBuT/Q+l5qOiBQoeqCfJlrBGIv5jv3RUs18WbZGP1lQLftGjaiw
GVF9iN6acKj6TDgtMr+2PNaJq+lUyVgGOCNXyx1UAHHt0c0LMX/825rEPS8yWKQPIrxoE8JxeGgH
nMZR9N6D513iEJbSLrK4UY1BWhGgvPt+tRGJ+GM51efOisq3Knny/Z6qSe8W4g1mPg1HePta1ID9
Dgm1HA5LQTI5S7RK9mxnJ3O5VrHlyi2yqeQSntIT/bjFajrvmICwhYfHpTICHfC9rJnRcxhFJBmc
fD2spm66sOgM49atJerM6v32/eu0YsaZwVckKSCt5d5KOpG/BPtTFy2EYFhRvRCYksl+8rTqIogL
/KLgXBWvdAS0aOaWY8YAJrnzFb9jNzk5MaGeCVuRD+rTIEh29bxOyrFAlmBhh328r4C+Lo1uHx3w
ZjXFGdfOq/0lcRkCJk9Sw84i/FSeK7pILQHlo0b7ShE5xyyLu1lzMS1Cyr5kEluaTCe5g609en7c
yCNgQBa+wnrnUUa9OqXCniz1UC7KNGYQG9jxeFs+pB+su8uct/oNkReF/9qP6l95HrI4l2zRoAsM
OYFdVjADaFgHDtnn1zwsb4/ZcIl5Q6Rc7/7HnXhuJ7vHIrBQ51gz5YgzZaka+RdBcdpYuhqju83/
n36FPyZeTQwJAyDkBcJzMdOjtO/XjMfRA7A6z6LIFgkMUBEPxNsupqxmzMySayel41ya3pIIcGGL
hXEJ3cdmMwljOcQhe2XWSne+cWYTBD9jdAMaFZZEPBp8hdT8OxSil2VdHoH+femym1jLVrNLPpN8
vBI0LfPMF+KTodnd5ZamIqxKfA4tAYpfMoLy46Vz2SRc6XEdMxW1NNVdGMvcED8U/7mGaV08hHOC
I0qAOQxUtvnWfIT9Wj90WB6HL8XCS7ns6Cz21i+ZGYJeQBFPpnR5x/l2e9Q6g95wj0Mm8juw7Z8b
Fhq0lYsZNCQ86XcOneWoKgPtEEhuxIIkU6JMVem0eUl+H5iSMBN+edy7Qeze2OggpvX65gPP4f/3
bFrzT1jOsQbQo2615VyPyCJ2xl/wjvSRSEr9k/StmuY5kZ5W0ANhEBy6w55RA24WFd+w2yAL/C1n
g23XFibN1iZUQffgezm15+Te6AK3GHXzSdk15VBwESCUTQcfzchzHxXTtNbnDI/kZYY7CaLMW4F6
QFQWjCZY38RwPOfgi9v4TdP1N7qcQ6DqHEf4KcT7AhNYEcUS34o/ss0gcG9Wj0pQmE34GNtcIPUL
Cq+PShd4zlB12oaf3+6xFcdjfy6Z0Yiz705k0SSIQf19bf0ST0BpHJTGWm7O75tITfPehZGf61EZ
xH3L1WKwkgOGCH4ygC5emsovwtBP23ADnsI9UtqnQv+vppUfdAnTOQNOrsNYFJYCUt5iMisauVrn
0Pb1dBG84xaY9AcceW7q3bnaecZrbCkNW0nHBBiMqDY+jnWCqCmeS7CcvlTj+pBePRO+6k2TrOIp
FNtJcPPDu2VjJT2/U64fgmLet8VAXkF2RwoNHQCWbyqIPK+v/pAOjYr6r2NXvTe4oZBDCzXO4DCW
hW2UJROu4dwsOliuryf+/KYlWK826Fn+8/4/r+6b53j/jMDUqrajV+bNPY+XpO6rHj5X+o1Yluuy
EgTgqYDVl9hqwifqFgcKitB8xv94T2WX2Nt5bOG37R4FmnfHwXKAWydkluE3p1d6hXkhL6t7VSZ/
fLAov3BivukUxlvG65IWkNSa/NU1VarVw0KZwo11zhKeknjZFqXFYMxOnxitEscfxPbIoLTDqsCT
eGFIJ19Zx1MxnZKZRalFOWCzIzH0vif19VB/2aLPGs35ku3uqCHvC7hOXLBdpeNad76Xm/5RZpoT
3qugDdvqGLLW4EWmAF+355KJuVGr8fFflrLmOl5L65HE/ScKsVMrK2cp4UP4Q47EXPkCFtmQl825
22/mwKnIy3iomAaMko8PA3Nsm7ZzD+yaW5VGaWDTvcDTz7U1dHZka61AI+zc9FUF55vq6cqBtjiL
kRG98VGsz0N0LOV6+ypHMoPNgiZgMbNPeWYcHpFbq/CvETRtgrpaTB61wqprVBqX6JOqnnHdy9ci
V9Z9w6plC+CipOtvhb/8NusMFtxaGA1dSKcsIDqmjS3wvZDF4+mof4kEjgzA1epLP/B2Bf+XENNA
vuKtRUPWgUwuwzzdrsqT1nRhQIwfsLodnGiYFLA4KKzpk/qQyil8lLb9bR6G2WLECBH3wP8IC4g9
nh+Wr+/3GtKhJwv1HC/P9fpKXf4pWuHmQv6jLtTwfgVImGxpvVt9jJeYQHSyKP6lyEXAxlEfpwce
3aS8+zJpQ4dqj8HI8RhxOU3hjIbt6mHwjKXzQQPhgZxVbcTVuvCgcol/rScvCLo/Xu7Hd6XVgk08
nW5kffq8YBkF87ZIyMYmmU939HTweoxvVKj8ZQHBDyIWPBLnqiaBtrdVqMtf9XL/0ID7JW+CW5xs
n3ojfAPYF4IWkg0f914wxrKqHhY7R8R0xflji9aQlo7Ka7fPwna/WbBlkjVPc+r9DFsji/zeRaSk
eocuaGPSHb8+9kj6319vMGDBol5SNJN5bE8u06RRSnwEUOOotjHaF/2XdqS8UUzIi2CQcYSAw5y9
2LKhj0g7zCGB0SnY1jptTVGmbMH9mzfPZ3voT73GxQrYeFq5c/fh4Xr6j492DTU9t7ozs4TcOVrm
4XIcyt+WzrHIuCg56YwAggmJE+0jVGLLX8v2G0pL2lAX3i3AOICXK6yZFuD4rAe903DJmHsydVMf
GFURn6KkSrVeTUQMnxWvfN/Gzi5keDj2amI7OwEiBUO7s1K9sS8PNlv/cj2SxvjiRgJpG57SRjh/
DxpSBXBUxTT2oQFIt/4C4XOrw0bi7a7yYNLmtIn2ctk+CpxsZX4Vz5Xh1LJDHHs0f0HnQxEgxxY1
wNptoqLHOAxvwBerH+uud+7pd6B0ptQQztLeXBGhZauWbZl0smXsguKtEFI0owzKGnfrjUIQZFCu
OYVI2RpXjunqeTmcZEKFZm6AtzH7xWa1Q34kP7pnFvscpOIwblu+nui4KgN3gcYo7sV31Cd+rFkv
Ng7Jfblj3FKxbiZbu+gvL0g7sXQeLjBIILrzEb6sgb2RMxlxTAWOLsQCkbg+qToU98HxBPZXPMAh
xXX/MuupXbOgPNxuSueKxC6EZbDxcZgIedcpaklH3swjLlrZLOfY8mRzL4pfE0IXXpgJn4c1q+0p
ai6tjjWIErj/LNWhYiyIjAn98rqt59ecMsV13tcS+SweQtI0ZtCXFwOMz+Ow5Vky+Jg0v0VcZkvM
cCbmnT9Q4cNo4TJpPyvyNArlSQMis62qREmTv7RxGGVcRQYCJA2Gk+vsZrYAY5w/m6fDA3LgD1bO
HeC1Jx6GRwNoGD8ACAKUgtdsDWcFe1rKyTY3JDPYjWb9UxkYwBcMWPLXA1uYt9S1FVnMJLgd0tEc
Pb5J/vk2tP2CZ2fh2O/ndYkMw6Y0Nea3EcPehNG1UKp2oxuvn2DIO4fni+2YuirEdBG/MF9sc3vt
Y2H7bBcBKid/oQvZUNJwWQzRsXVryYNTCnjkhpYFj4Sn74JDJKRRnfcj7jQAFX4U0ET0iTH0IK+d
oJ7VGy5cx8YZ4aGHz+QuUJ+3M8nLACYQeHnDSDrs4GvLN0qrmcNGqWb5t8ADvzoee9dc0dVMMEBP
qRR+vHEhjV79x0JpjLa69WgwAF4rnEBw+dH/HoTqguuww4JTvLs84CR/+zY/vTvrlC/VJVR1qiOR
1I1SUFeU344NnW046ZBqAZLY+WGmIBhW0hqLc42uCaZVjIMfBPUdl8gJ6aagb5rAzZvyPoF6nrqH
2RSorUzNJgkSwMScjv8ZKAtt/OjkvTt0EQZLEOw/WX2p/YqlUmvlKirN8+gyGpYLZbDZyBLxmCW4
+Q0+83hJkX0I84VGWLE7aSxISbtXIrr4E9SoRTsTUUEtq8e1JTacf1UpxP8Z3hUFOWUYo3J0d30K
EKy63RNFfKzqYeTkLoxwPcwvkH9SmYbsxR/Qs+viWp0XwxLjWfDcBcAfpwH+2/ZzjldPKn5ibJY9
40hCsnH7yJOIM4ad/qk9Ksk0T3uHdHEWftuYR2r+rDatDUv2oQ17zYHXh23VSMXh5z7exAcqvVrv
v7ZYI398vN0AKwePUar/rzpVZ3oBSaZWx37q6tu7m+L8KB1uGxG61ubzA6TuyJ4kDaCzvmutEOpz
2VpTew6ubz0GVpuFXZrlcpKxg3b8raWDFfvMfhXMrQ0HLUr1Xu+5UfTnS1GIwtJLBkQyXW72iuR8
snK7US63HTOTc8SRxwDgLwSKQIDww7KEFHVyakeqoM+2bzQQNPcZt4i3aqYioCGuzneemE1pnBaD
NgHzU+sA8mkymAVeBfuCRrwlNp8BktBPHUTyFxZi/sPHomA6QsN6GZu18KXL0bk+jfinatVSoUJv
ItaDCZX0jUOspj6mCTFEzFRTRz5470IOF81AtO0pZ3xYks/ptbVZpVw/XCOtVW2hLSQ92UTLTOfg
Il12MY59C4sy+a0R38KFvgy/sZH3d635zNZN7Qgkd9eQDQ9YPYcTPzihZcrtn262iLGX6O41va9T
n519kk+Dy7UjDKV7gaiwW3mTCYGTCCckNch8yPmxfGnvqwBYHP+XCUs6VsbukdlKvaJAF6PsZxXO
Ra8/aXvH6PSaa9Y2tXIwhVW+VucvV27RYqEfmT2lHZ3xsA+L3HOpI0tzRxt1IdK9+TTri9ypGly8
oJj3MiYWQZGeP+6omvkTRDChkHU4xg4fThqUs7eTKQFcDumvYj7aCwA96ZnkXyY+zap13nUJnsB7
QkN6L21POAvooX2IXLUyD2JbeKTwKKXXmACJp4oWhmgCtCjq4VQd/kXZ0XEaO2xJeUi5ynAPK9lu
OwZP354yLDKO7Nb/V7rFC1AFDKwNbo8dTbbIf7HPFjEFDdbT0qPU6WmRZ480uPc1WNbZ+pRu+vvQ
cH+y945XwLr/MAKRXD9F4VzjfBnkuO7NeBPqu8TG3/XEYE/vdKt+BfHrWd/qp6umjbtNpJditdkp
r6ytVaZL3VjrwYLQuIZwAFuF3v4qYz70LkC6ap2lSjc6v4wDFEjrwditylwXg/hli73HnmAR+0aJ
f3p7mdDJJeVguvBECroJG43KO6rEIp1/RfKczf4orQPvxocOIP5HJmCFmiNgSxElo6rX6klNDsDU
ZpApLQ4x26HrvoGoqe8UHZ1qDQVqK95scPic3oxKUkq4likcbJfU0dizsC70eyQCOoKrQB9VMatW
4qTrr7JBbHmcQrLa32y/gN5uGICtLJvfK7fMQf2o9RkROBiCVqJhZDVRay9oAazXNNcaKHTQTlpm
DgDTh7xmngQSwuTWrppsuX38SUieXeIp1QIv8M4FI/JLmImMUt5JcBWTqLuM0xrR6zAHdozWirkK
vdhNQ+Pto5munlunj58WmraLhNxsV55lHucNLXha40OFjSc4ux1XNIsaHwm9kKQHaXpxtDYBFx4j
ffYscI8WpCg4BSIQBqpAR4JyzO8oVSxU1RFLhLL+lKLe5a9bicbJYKcWacIgVosf7yg0O1bgH5d0
9Y7URYUMkf3nrAB0B6VPk7PYVmD0lH49V/3QvgMDWnG8lu3g4udqmgfJUkpHjtjL/+z0zVXLO2nl
4PcBZ0NMJymkAjZDc7JjF51jscCtcY6/uv7digD896UROvXvwWjxzRdBwAZI1aSEnEQVTn6wAMos
+df8e4xjGVmsAfak9djKwakI3RdbhQFsCxCk9aa/K83iEZIpN0jbdmlkAdx31HKBfsjzfg2GXyP+
/p2C0lTVlB1+ge33qNjkS3zbUpF6mnafXc8ZDtRmsjKs/AKWjTbSakFYAVaPfaS+1Nfb9oX39kJQ
qsM+TraHXQjpu3AKmqv6Med1xrFULYRsxX8gkftBXKQBQdORIfOWFexCuZGp8elNFj+osm8H2d9D
8C5WGiB8B0MYPidf/P7oSQ5+k/NRz3MsGLCSV2dFT3fSQ8v7cp++qzLTniKNqKlhRw2+Hx8nkxFc
9J96DsFNgc1kvFbGxsXKyCGSsI0YAsAmknmmwY8estPG7zqMOcQZjRPBzaJ3byHfOFNAi4UhqA4m
v/J1z8E/wC4ZDw3S8Cg5M7tHkPt7rdPaoHckAalFVpPawDBQP2FW8vHDuJwtcXyJdpHOwri6l44D
3oQRC9SwhCiVZCFiMRqwnz1oWSK89w58+n1nWrzOD5smO7ib2QrmMkZ2d7SSL0dzhrIczhx7aX+A
9d9K8KFLqdFNeq1eqo78ctbRuWQmnA5aSOvZwljCSjJwLMmhDf4a9Q1ObGLFIlqIXLOKmyVrAdAP
QFneWCLp2l2+4SnEdV7iwQusc4L7xCRvmOK/kBBjhFFqrcKHKBleYjpdGr5KVqH4ddwyShlUoaEN
cd5m0+oCAaOsIwH1sQewVRr1gtPUsu+JyYIpxIjVMwI/CYVpSAKARKZh0knt98xzKYYj6t3DgSgw
76qkLcTgCSiUofNz7PlZyC/oWphyTQrfzKlmY4CcuNG5fO0k5Vkw9DTVawrO34xbtVHNtbRes6yo
xSCexOw+mePZ1FPijwcEUN0aTEP2H4q/njTHhcnXWmwXdgwS8HndQKYjVXoHoU8/R5F53Py9rwOJ
XfHg7Z0pD/bPUZbiBbqQJcSbSEJYHomOcC1gVXYLJal2vYk8o4KJRtwR2lV/OCOY09tliRk4+JqZ
kv/S9s+CazJpT6tyQ0UeYMhLp3XR33kd38kwCRm0XUAGIWPPgg1BPkJTi/U4moNVk8JAPYaFrud8
U9+4C82hK92uousRlS1NShu0OVk5753gtDKp0Nd4UYRTMIjWtT+KqvHEbBXnYwaEDZbFRQbXv4+Q
BtUUHaoWh3wk6BdFbF5rWaPHjeow1L7OgHPzkjfnS4g8klI07hq0DHC/wjMvXFKl48C5p4SNZM6e
xobhPJqFqKDCpjhSrgbo/8AtcugEu7qoZObnOEKnhFMSoAdCBNg3k7xNWy1muH0tsFkGEJKmUNYW
sUkfYqh2HBNaYM5m03uRdoGbLO27lWUBdzJgJ/sn5DqJ+gF7Ds5LIcUsRndP2P1MwgeJ3ReFVUMK
3HTiP/EbYMltfSVJs2VW13LOUwpouq0JenqAPa9t+uQyxVnIOmBwOI4cl+A7mLswur/MY1kaxWTK
vFQVkQ1G2RdpVskRu56wjWGkmBr5YAl7EJy3qv+HZQGCbmYLWh+i9xIplZUnf/0dhnvmbw/sMa4O
5AoeanvA6RyYHDVkrj1Gg4FqCqktb0GY59ZruCJCUpsVPAe6xhMtnDKzZYtejJv6xWDGw8qlOBdG
Mb4YFFyiWVnoyySrsShC95MFGkduhN0tH+1A3EupfeNBePIprRtdr9+t8/3+HRlYmG5aYSqx7S/B
ooqlep+07cPe0tYubRxGJxmH4I+aEQb6Qe249o99bSY9kLYxtkfBCGI6wfc39acZROXd52qnSHr5
qh8snGdfD7GqX8BspPd662W7tH6xJ5mcsERCYpOiLJuW6TBdhKg2PUT/NZwVciFkb/3uH7MqPh4Z
DNabKRN9bVK23gkFb94UWyDEx0t7EyEC07YzJl62CvKf5Ip1+8Al9CVxG4x3uuIiKLaC/wDRxuDa
jycL1bmjRNCUhIwNPhCFudEq1YwmyZJ4TkCzG8iMKb6s3hSZJLvlSSatAIy7//uQIFgJK3teJI95
puVwA9cf0ZDG5m7gMTH9G1M17dmURevlsCeAtSQ9SDH3It8aBUNoNxqRPWBkCJV+iNTtcJraQ8g7
4DlqcumHH+uSqVkuK5z85CK9LT4cVuymEH7JGES44BIV+UuzfE7pkIUdaAlLD8kxxCkYdpYlluEz
7Gu6dY/YZ0TTmiEBtaP0qmmnjZoJYVLNoIVEzZ9y5DE+/vZP8VZcGD0ewzjEiu4HpSxohVzLyCxK
4cNczJVmbZ8SOyCb9vLPK/nl12igIA+ObkW8RuegYtI19YRV3iTCKkiCQxH5e+IyBvTR+6KVrXhT
VEq8TQYOAgIBqwDBGBC9iNvxZ33GqATX++z/BaphUv8cmmTn0Dprd+j3HFKtkQ+50heiBQD/UhDq
TdJsdSMppM+dAy76lTGvOhxU346A63IKIQJJbgAjKdBF+rEMjNlgu3Un0TCJ7BkqTVdm3tsOIePE
x2W8DI613FZ5QaosmFqDVdoyj4gCx/ObwExBBE/s2Yn1BtYv3FaZj5MBp1k4TLxusV5TbC9+V6P+
dYMqb24OoNTqnRWpKECFJMEdyO3EZ+X8uGid8Huvj87tUJxsGxwG7wiaPT9QmSm9UYqpp8UPqd6q
gMuccWof+WUxbOHDN6/ZQU0TX5Zclc2PSvBXydqQhaP6fUOrRVouMVCroRFtQY+NRz+sonbM86rB
Cp3eVx3naLL6TisLELHVbQrAhRpxYSm4lky3XpIGcfrcIGQdAn3/eu3+ZM+UtGfprSDIj9QoLdVi
I1M2H7NgNKVTF24Xpj4eGRtgDzzy5d7bsvUnTvZheBy/RVFUNkCLOGubFQJxyckfiJrg36RkZn81
y9ZoSLYTLDRGH0zN1LGKswgV3tBSepvHavZ0n6TgcJ0csEBRN8qxnzneM0zUpyjt8GZL0IE11VK9
TbY8Ws06RUJP+dSL+t3G+peS9cenHeN/zzPluMvaywPyve2hYyjtCRDWXNseVr9Gm6JAEezBl8v0
R079uLywUQRksGwKXd9dgdRbxNfj7ohCA5eV8MuhEmKJGqovYQ0xcdAO0JUUEq3RmvErWKOlcN1E
IFuVmu8//XSxcoObNDypiVqetBYFuj2289vKHXDj46EYdiMM434SW9YePjcmmQ14bfAjBUQcvV33
dkr2tmC1Oy1QxD7YrJSW2FPcAskykAotA8n1LPTCzsnMylNUVo7gfBfI8RBw+naQkFmCurX7TF0T
uVv4eqgN2pyr2xDeCt/b0XJ/EKQgETt7op172wtCnInES8Fhn4hMrEDognTqpu2q9Q9bxfmPQ0YI
u6xzPjfmQOzlGQMC5Or5VrvyczgJQBjfb2YDW8zXbiAc9PeBiF3HcOe/zxIkXVgZyn5E3davzgv8
bvB3DVboZzGr628EEhDbi2i4+oB0S3d/m0vFKDlshA6TiTsBF0bcKonniw/1Xonke3reBJwXkaau
Ep5HxHfkW1/6AETbGbEJiMIEywbatoxMADhL+yz9UrBUqPDOjAWu3baMavgK00mIZLV9lczjcTWj
MgE6ugSnchKQ4kYBkDa8V7WQIQS3jS/n3C+83mk7P9HfX60F6A5AC8ZXkCKJcI3mvyPA0TuCbst5
RFToDwXJ9+LzA/kUpY/URJ0zLeeLMEPMUqOZZvjsDxZUh1yI5RsojpFpnxm8GCLiNXjW4fwDgLN3
R7nND+kQh5H7uB6hSfLSOCBurMqwRzFDfThBPVrXJTj7QeQHnm9JSLRfpom+zFgQ4Xw7rSclhi6S
jT59pUvE0d5oteOO5V9qAcjkLB1kOV/Zlmxy3Un1VzZ+6/vDN5yEPPyQzopZ6ZIwzKV6e0sxVA96
qW2XuDyuGWVbfJbUpqriFAjbTyxYeLvgy2U1RGHwk1jdK+QqWNhNIIH0s01JxTGth9QpjKBpx5fY
5pwC4CxCzV39VJnx/EOTVRXLX8ELe0j/dQ50aI/kBVvq6GbxpwQvYhIONVJCJO6JraAMJ7uwfige
3Wd8zq3u0BKhQ4M/1hR3j8B+h0ugR01vLUIlQ6/Wr926YW5zmmjYSkcdHQLQlWU9xVYwfeY0YhRQ
UBRbNkgv54F8BfCB48qeE2PNHSF/tjLFEr8nIekrlwn0nlM0IU0l3IESgkiJG0YrEKCTkeunJ0bU
wqKjL6++vKl3Cig1YKA+KSaCxOVhvc6OpZzS9euX222j35Ow+fTVpEoxPMbKSmvcPQ2qKOMq9/kO
FUcWQ2RNThgc7MoTa/LgO+orECXRLWWkM6IUIgrceDD5GBwbUbR9okCOacu+cD5+jqd5a8gJbhkB
G1kT2BPENvWlUQ4b4G1uKqq4i5D/Vt5Zp+lylPoBgFFb8UrKPm06q66lrQWmlRPoEabZhC3cta5t
SvwpV8wCNC+QuLV+1sb3kfqg7zQ0L5xLYric5hANtY47Q4c3nahZH/ckHW0W8VGfUMGMo/vCubIX
SisQ/jMOch70Zb+XbTB269jkpe51Z1jWexFGHqtMJL91yt2HiOeYf6l+pnfQANJZoy28BwmAkv62
a/Afh+X2eKRCYo9kN8/hDXRE5fuaPqgWfb9//8DqmL5IVzS/PZWzKE6h6naO3rERD208rO3TP7Il
F3/Q3aJLZSLfRjOGmVrMu8ZNeYDzfGQ5EHv7qUSyp4zdQi0Y4iis19g1zETX/t0F4F/7GHPKwL3X
hUKj9+b5rSJgC+D6YzHlNGXSqSBeSn3NFUFBuhgozaLDz9EnrKlrvE7iikXzk1UpHdp3Smt8Ztcx
WqfzqK9nxdPyuwd3ggDCd+FlC2K/hvLC9UQWnxrEmf5itnNF/4oK+FhUJLOm/bElwMtp/RdXT+Ge
SEwuzrczWQ+VZYnAzkSED9i1uN8zTSoS3knTdBZDE8CUUfCW1XLsLSaKIm3//9a3jBj2gwSRr4H2
Ctq1OyL9laeu7QI01PuVXTo0FwFW3K6x72TnHScl8oCcSGmw7N6OE25zoc6RqHgLZDV5mjaolW8E
VIwirSFDvqdCMMlD2te4LiBIGUO2cTjcovf4nsyLmE4laRmZs2oJNqCJeljGE1EGwHCr7F5PHNAf
aAzkzn2iI6Ps+YETiLwP8P7gOD9bIAtluxPkvQQT+i+HIrnX14mJgA3HuM6VYURvhJvYm44a4b6U
WtuMUtvyVzoT972j8Slwb8nmVakOzOdsHgcaU0nn64d5OC5jAiwwFtLMJEI52PtMwzxqjlCo5pLn
rXMTnnOIVR4h31W+YvqhIlgw+kHfPo5+5BVFdnK0uYXQha0uhd/YpIQFNvYC9s58wopDDR+A0TQF
lrpG8oW4s1RqPSLlofKh4TiKgkWCgPIO7NZ/Xszhtntp8nR5ieI9rhyTU7khu/5TjIeYhCX4Y7ND
hHUbsOFGxpXlyfoq8CB0IH1IzAGAQfGVcYrcfvP8cWEJKMy/nRUlnhq99/YTKM0AOm/7cy0pKyCS
1CnDySVb7xfsmw6TmMoJ4Z2RAo/7du3fru0tLJSqn07xYBsTM6qXE4dKH/LhoypkzbNKuUp8wacL
D+ADzHuVlDNzxWm9SMRA6Kk3qiBvSHq7TSc5qUxl1d4JOjhUY6jplyeIz0BjWfohj31v7URr0nD/
sfkUhZTDP221Mifzmxq1vEmjNDmuYek7DmqP0FZi4rYUtnRXxYpH0uZnVdVGplqWLMJP4bq8TqZz
H7DiMz7xUhIaB5SQEuHD0KJzB9fo5Zw2OmBcuPvmvpunkL8jxhWL3hNiZYuW4aHJbXJVYgc07xGK
T3i2K1174fTNMDJb8A6QB5ngFxbotQ4wbKSUMrUg1S16CyqOEC/A+ftzUuZeA3VKfwv3Z7WsdOvv
zlww/psAIiIzXT7iEAYj05JY/ey2Sr9xx4hW2w8L+0tovtsA6BGVsd275GSwfdIu9EdMKSdAMKIJ
09MsUv3kxgw1hITXmWlt/qlpgiectA0rb5uaDfGLkXTQ2HZwvXoQmJbyXpgNyeIaDhugWj3rCdKo
EP1krLnuaq3DMwKZirGmMHIBqaA0sHNcnH/yStlPD40PyrXtLOL9ZtKVoM3KH2ti2jDs881biNsf
yvlShSUyyTatx3Ex1ikk2Ac6oJFYgZV/XIfceZanjptyKQMarUUsbN6zvfQvNJsrZPu7o/tNFFbG
i58Xcqcpl3yzAczKZY3iNBOTMkjJ2JEDN+R7uM1G+TsYHVqMtR8czm4R7YkGBEOMi2ComwkMKOn/
8unclL4H0hkkr/NLXqzb0WG8rJgFIXxWodEZXm5Dynq0gENApeiBErxkxpgi0BMI4kla1QQHkTLH
W2rOuEfFbvIjnAO9qDtbxh4HcEZDpMJAAoXp3YDgNg1xc3UlGHhaZpZ5SF6GhYtYEfjtBZqpz8Jr
sAV2bsWrWXl2CACB2jjCPr9fMKBlOAnG7mEhty55h5zwo9q0vZD+7PPqBLzmsW3B+x6g4v3ymPeN
sZSU/eCRSZ5DJJZ8cW+FHf5wWOSIq2y8uAoIbQqYDay1foMJroMesWgcUNWkD/VmteKmjbiZMuNs
33kYK8Za06S3rSZhQH4IjamLFtMChBkgYxoM46lQRWOZVKARJP70Cn38W+G7IDzBI98RleAbJZxp
UnZvuG0eyUb5WdLeW0bsQ1Bn53BeZWVufIa1S0p/yutFZ0Fak6g55JBq5Va+EfXeXSnIbT3HEf6V
4SW56tCbAK6vYd9JlQdgZHIgl/h9yqfe1KC/6wYdNKbaHniiCRJY7ocXW61aLHgfp7vvETuqIG7x
uj+4Sh0U40djsX5eP8yiygRRu0bFDbTRPhkBN/6yTqYuOc6OZp7lgvYYtojmoN+2TNhaag+nq4WC
IgMqGtDqSjOZeyoixpgFqkMGYwqIEIDcUa8iem+aWs+rWRJG5sNLkTwZ8lGAIDgdaTcTspsyWpHT
DId9TBcwg6sKJ0AGsJ5wgr1dvqLs9s6Lm9p88d08/KXwsfifCFXTtuU5Eyg/0274FTBNUmc1Zo1B
YcKE5kFGtthmXaEApxrGosSr7OQ2YJBmYsLPYOgxeHz/b9tQkS6Hlu9XMLqhRJLbBEhB5egdkaXz
wh5v6VNZv5pf2B1ixD8CpR2GGWCKFRSWdCr6A6S3lYlmNSy4YuISct/kMDKnwk1lpgb4paN3DDFD
OHgYi4sPVvC8J4FyGO4OcgASkf1mdmjM7s0SozyV9fzXhfRDVJ0smImy+Br8Gdenls+vvogiw7fW
+G08FgC1oTn+l1A+DYe65PPCQ6vgj2UjB285GB+PAJwlnlpHeU8WR4r7MxCx/1S2gahCtYkk7Bg0
UJeNbMNbfwmW4n6fyjIKNzPfibFB2oHhIbX1YWisiqjfhBLigXB74yPfjbhsHyE6dC0vfw1NnQqj
WEW9TZXDup0XWUplw2QNH4OCzZH7qnm2SCPcNTmdJxj+XsyoYwXeVdmX3LxyyPa17t7jIrhsVz6T
q9f6YTtz59NF7/ikGEZomPVleZxlOzJfF1s326PuLpbkWq+dZVxSMu3ZrF9oljLyo+oRQekc18pH
qWZylkfsxXkqLkF/klLJSX+GxlSsJ75H/5SmLwU6geJZaOD4ap5M/x3s2K6xWXOLwl9288TjTPWy
s4lEb7JbnmcyDowJLUXyWdRrXqoOCiv8wUGIYMR+nkRBqU1x8m/nY5zH9oOwBPldu558IaZimlhF
kbjHlLQVrEeC7etQG/TBa/HtGw3CXpgRR4nI/dC0eLvyUVMhYvYv6Tgj1DEy9Mw1q3b62ygYUN53
/v4jzRqdVr0VarpyOtbY9UevClrJps0jCUuFDXrH8K1yt6U0Bu6PrqOQGjfGA1HLzmZE1PU+5zxj
mJ/mbL0rmbOjliaZC6/x1JBz3TJL7CQvotR2gvXfMA4rltGjmvRrV94vGHpy23V0PrBdLT2ONdHc
xGbxMkHhTohrs30cDOXxIda2+qth1m0YzK8wtVAAZDtLoqmCA886WmphC0ZBpau34JVPFGCYv0EF
Xr6NGw/Uk/DMns0aVrqNV2Je5cdKd3QFsYf3OeRJK2sH4/OhMUyMFUdHkJtrLfzxkV+u4RNh2syT
sR70szZEOJ16NhkX0TEpA+Uu9PI9DRXbM2R0p5ewmRiG8zkgJ18nSNPHGUxc10klRm48W5JQoZPZ
Hm5jgs/chrz1oMdw6Y2hs8L0cV8WrRf1lLCIAoM6+taNiNFr4qux7mA8wkqkdC0QldTDheSMWfmE
45VD93Lo+pIehuW7OvN5hFBvRONb15g+Rmelg1srxoOO7aA4OBgdfUJ4hkQwULrLQ+eXvH0fpu/L
IY9Rk0VDL5xmjwhD5Sn0KtrkV+BI02bDy9jdkvPlJ90DME20+M8fqLQ179uV7LbnsrPoF7SgreUD
feVfgs/VbaYhXA6Bd+BaeJTtAzM9fp9BDsxFpCyaEjEH14pJ0bgaEdiFuUGxNW3OwtA3XenNOqfy
jio1SpzCjP8M8jnVa1Oge+xtnK5KPOJD9jrx3fHlTZDS0sFLxSvIxqbhTNZ4TJIfUHCf6Dl3FGMG
k5+EJg0Tg2i/7e1/GSSgTbSIV5mPhb/4ZjzprEBRVauvgq4J9hNi/MKjn0Fa24lYwwS1Y7z0EOKS
e7rB1Dk583FNDoH0eCdPvYDQbj92D0/z6iHLh47UadPyVEYMtwfPH7jpHHP0V6OGxaviNKeC7cJk
eAz4a9h2oIBbqqPlj4/i6skvTHgp71BMHiY8+o/RDsYWkOdIU6z3hZWnWLkYDrWNhJ+vrBAlT68f
fKtVjjtd8f/GZifxbYrTG6vHxXIGRzxSBMBFbYJEfQDdmqS7kNZuv6Sj9T9UWUuHC2DUJoodahyC
3kir6ucjSHptM+57vxpFpr7HERwwfOsgouVaPBaZBtFun0yMiBE/blJNdzbMHvmdTKKWeqBeZEhC
isP5RqDohathkPOdKEzK8CePzh5OMLL1fUSgAh9Y2IY/DUFipqxgfheYeIy2s5ofpSr1kqTWxbE2
vAVJ6PK2MIaU403AyFg8NS8KqXOeWXzFhXDcSDXVB34OWeiYbFixSZ473vRAQxxx6BfLYgczjmQs
OEuckoc9VJN890+zZr81eabeq8D4TbFYoxuWRZGh8GOzFsxvtOlpww4UpGsNH/Jvp9T7s97jeuNU
ApCK4LVi7VbmlfgoyoHOjbVFOWhJ2WRwVJ1ZZS8wyTdk6RpW0TrAp8Uh14jUYEZqT76fflqHQnn0
sHgRJtCWY8/dvhtEV7LTd5Yxnxt8R8cWnxkDsxdSB+flJqGcVxWO3aTIdeWZS9DFHG0HxNhDXT69
CwHChXe09FfxyZroiqwirarOp1cQEPuYivHNA1aAw14OTtP/UVQ8DPZKvhQtQsm9tC+7aH591sao
ZxSMxodeVnAMox5l2ldoxJ6Zpa3pq8LiRfCr5BKhwhwWTjmMCCTxq/kuPNOds4nh+Xn8KXCGwKVI
B1rNNyRvLlIA13Qdq2BNWpfhsuReUXZiG+9itWxtS4suFUqmKySAZr+53kdp9as3/q5CrRbmuWJI
LDtDRGUNy1o6l0rhIWOYkFAkqBlAEKMscw8ojUvbgVxUBzdhqFQJa6U53UrHlMmHYIysNzTnIhDJ
T9Mxspqs9SmnEmrhV/R+2FIaGDYnJu/q6nOo+4oIm9qRjKvLIPQdJruWyF2JqxATh/RCWQzxIUkO
QzrX9CdoNF3IFsKY0aQU+IfTaPNwEY5yOjKOqC3mTVGP022Iew/ZnFlriB1ZbTG5hhiu7UsT2Cth
o7kW0Nb2Q2ZVRyjNWoZX0Qceu69XwXO//3ln79LynZEWJHiAKucO4hsMdnpbTsCFpTLA25IFZxGC
sJJk2/inAWiG6rFHy9mcBB2zrqc3WxV3g4DbhvUL1zuNwH+DZLeYbjweRdZ3Q6Lm0sbv8bBsmxWo
weP1O6zMmeZuQj7JuEkWOsOmjP+9cxyqai663tz2DUGGZgFp0OcTxhfEFQRIuCys6Vb9whKxy2pr
6GZe1VMcUXi263g/CyhkK5ikqHXHuujDHEYamRYO8OAslv83Bq8Z5D/2nOjIZQE5l80G783h6pBD
4aaA7vxE9T1hfAg+vDazGpynOa8tTGGbjc6cTq94IWwXrlRlBIKAeXXUfXXmPtMB+FmjRaifDziU
W1puWq4CV63rKx9aEdpMGf5bnfZwXZ04EbC3ubzMrmWJqiTErH8PLlh0OC0TCV+Ew+h+92+AStwP
tY/x7V0o+Qqsx0zDBk9c0XGdl+NoOl+Gb4ruEVJ/3lniFxBJ6GA3vSIryl+VSMW7hGYmDaFCG/YS
N/ELqmgvmRaKiEIhLg9eG8tssO5/QmPihC7wgp4ghp10GS47wAy7ffe7zMY0n9nN/osxdF1FnUKc
6U9FWDdRQ+WsCMMGqHPd4IItcNv3ZLlNVNX3hY01Z4ZluGzDUSyNhk70Y3bD8AaNi1JMjqXs2AJG
sN1bKtwr3PmRZ06ySvVvAcDZjTovnNcYPqBC+B5si/IdTaesT7RS9NOGAAqRm2xboDNx8AuMNtnG
wpn85Bv3ZDQiMlweOzrrVBq4xvo9i8fAkMwm4upuC2Ry0YPquuspPYLAEedq1NNiDUrjiJv45w/V
7WTiHs0VTGuGUcDpciwP9OJiKlBMHzJFNlAoQjuXV5nUTh6nYjerNrr+NizrMB4QpCB3WOhY5xoA
n2i/H12iTEArxmurKeZ2dhEsKqUWVZEAIl7TmdFX8VrQgKh7DadsNpkSavJZtEpnsV5WAp+CClu/
fIPNf85r/q3o6k7r4Ml+NabecsNOW9w2iDy6+Ym3p8b60PPSaQRZfzA5uyDWRLQuVRZ5rqTgX3bv
bjKkFwhERkznOk+VPyLsSzSwmorKmBbZUwlwkPg0Ae3idqzycv/ucKM9xAtSR67A71eEMvjAM2BP
6yUBivfVsGLy5YHD4CbHdiLL8ekrei7XJzT8U84MtPjgPmCwF7xtqI53VpUyrRBvAFP+qMRdIA7s
MZqIggOAYuHqYundvmqLxGQmd2DhavT1GxvwtQ9+5qUWvplnSLwHqzPWU2wdenWL3l9iKc6fyT2i
q7Fn56FN26oQL2nlHB0EWvP1i6ynUtg0tH3/Nk5sPJG5EY5q9lVnlUqjD0Lj8U+D9fFbvxJRhGju
FmOj+k8Ab/CHAxOsnojjOxV0nCvedRbm6zM0fPTtpASB0aqFq/YBiyU8D5ozTkQ15PVZRgVhdord
hx23zxflNc0m9P38kHxKv1OQ0bK/kaB8f7dpbvgN6MBXhRwkjLZvZVYsTl0l+bZf6KPTUA+zLlFZ
j6ct232eX2QYgnTLTaOqku8iIjiVHItZyczLzl7G/SeEkDsN1VYdLRVVunO1XFm5QyJmoyKP23T/
p1alp8IRkNOhx/Z8sK2KjnHV4YnDYhf8Da5fBV9Mt8YvpQvkYxy6C4+porkOvC3zgm3QN2WB/8Ja
249n8t52jFOJz+a94WqL9GAaH+J9X8kARsOnzpZz8Q40MoeLUvknv1y3tA30U0tdGaPEcVV4zevr
qHnXso5aSyoQOH6lfPTdKqx7KUpN/HOVV6oG/n8cM3VxJmxWZpBrKEE7Nydcfr9k57J5ZN+ZVdWH
8puXNg0fXLFSgmmpDQq6fmaXgoQrGDoDqWqyZ7fC55HRX9iE5DdhsvIAYew4VXVeHJ3QhKZsmdos
StlatSRi8DXnez6KqxSXGAU60okvzFp7PBVNXy9EG3teVPWh0Q9c5lPcXW0unD+NknQAyZwacc5y
xa1hEFkWWKIAtTeMExiEfIR9vCJNK04PYkk5/aOzbRB33hE4UDSblpuOIj1onj6yJZaSkfC4u+cn
Fy2Es8WfMo/9KwIqJIin/F7viM2D7LSHxjsm4LtGB8WKHdMrLPE2Jg9TqvIE0hzlB0NyvR3Sp5pe
o+97KAdDZnnIshlQDwQixARFCcwfXdaoC+5xuZRJfmXvCfcb3s4iolwWkRq1mWKA23fKHMPwE9BU
A0pXhycnQHD2Xnvy8nLPwQo26OHrJTRhlg4a2nX3jVsGPlHpF8tthGCHG4LZiV6iJgGFlIteq/Rr
WTpqsX8GvE9FOv4K3kfd9AxPBaSqhTdSSYa6sGKOWaVp4OegHKG7P2tvtcqEp2GuXDfQHOaeA1aZ
n+MfN3sba+8dibEpczQqAvDSQomc67h3lsZBBENueQ3OyPlchrnXtcDd2KqtgCQiRFGo/ik1VyDR
EzHsIsd9Hjmhg5TfbvowSdA1zC0FCVn5NFYteOQKw6065lRvq0XCtg40dnc0I/LVb+pNN9QHgjYO
Jeqq7akPy0zLv8JCQZwLlZBPnLSJL7POqs6/A8g/ITsSVVhDUZ0VdylMpGzB0uo0PGXTtwXPjOa9
vwiibqEJIkkS4U0XqK2MIU52h7i+psohHtb0fEJ9irDcw1nylifuO12C2mCzUGbIqhz3B4rknsHc
h9LVQ/x3qjbz+Js90zlKCbhvm6SphumfzxtK+NNt+rLb9GfXiiV4vo3qQbQG6svlMI71n3vpV8Q5
fjdiMZki43/86F7VzOmqof6PQodcS+hY2iyloZu1OA0DkJ6TgMXQq9b8OLsbqlPTzH4U9ywe8Mnq
eRxe29/VH5CxU2WhTDM867a1H5FmcIrM6fa9hwcf/dMKS+T9ZELdiY7ZReN/fA58XEssIHyNBpKS
KMzTxQS63LCD1ftvG01se2yKbpZ9tB9ah0C6csJLLp5e/fDSctB2ZvtXqv0/5Vy+ATb3K73iS5JD
uQsEXuLElu79KpopN4o5Wzivxlf2ICQRJdXzkECFJuMIVlJ6jvoIp3B752rXa1HR8b4flmt+jX5O
TVyXRO3EezeITrDQjJY3PjUOYRnWAQUQxILCEphCzlOkohfNiGArqaKaVFIObANxPYSRigW3CfLD
cYQ49sNFfjhKGlyzloKh99OC3kRX6vgh0MWZY41tz1CHXIi08nNvOhzWODADfCGmxlkrOgAESIdP
i5q42eflgJT8x9ZU/o8p05+26nB7u1hpuGKYXy2nWvVo8mB6DcOHEeoV2R6uW4gN7On9rwayDAoR
yHkFqz8B9GoLB5gEeJ06/vbpq+5rdshHWTn/IgVsI7OtM9hfyNF4yxhCDg5YWw9fwoUMvpnZxOxC
I0Ew7XmKa29gCaFMr7eGfnX5uVhwjjatjfe8WA8GkCiApGt8F4Hs9eCCf34Wp1tFJt+N+ehCyTra
W2qJU4XbTm2zbCUEC68QkkYpmcP8dpoXQOsq5x3cwmnQ1vrwtysE+xfu5lPxfoHuNf7OGEuQEuUy
2zw1JN259BS5Wf0G39B8R6W3lb2ElJ8t5LG9d3dSocQIH+/CKstPOvXKE+fJh+wDfXW1uc8ltO+1
r8/HPkQDio4pkvTM5OVv8YWnU7fOt7zRKkBkLEk7Xl0CG8jmox1r9Yn3mGatIvpoGTKHFlX1axHx
Rg4s9l8H7wcuWV0KadFiRXmIChyKVAeN0s0vNb7+5JTv/+eNVQcMYfu1qstwdHy9RHiwXPz4P1Zd
n68yb99xi61ISXcGmC7fq9DGpQwR7EB+F2U+rsbi1IjvQUCsn4VZpAuonAE4nRq9Yx8iodk5RlA6
MovpsGH95YrR1B2Du+LUpbMUD9j+rXloL924eBrIogSTrpwGhMPJ5wSJtGAc8iGOlBT0rB68Wn8Y
suZKB0+qNS5E6L6Nv/OFKgyME5MW7tKe92CDnigDjKjDElTk/Vf4gPlqNaEtuFyGoBPeFWms4Wh+
KOtB1hO6yKRWJTnBwJ3V9Hd38XkfKAXpu7sUpPDu7eXrnDzaJ29jd6u9U8mkyvkXaIwEgFfyyGOV
Cd8BxkYJC0mjyoU9pQgWVz9nm8aDu4iNX8iyvSZd7tJXiSIvyLZkMPr3Q3034yYEuf4LZUmzrZ1Y
1TCCYDw6MdTthrhxAebuGa/wGocy727Lof4PtZDt2EJyvwVyO6rEO1yLHkhrn5lDFISQXWhbtCJ4
HakP9lyGAUpGROs7Cod8Jb/fiu3ynkzfp2LKk/nI6lYN9UlbaWpwi1BqPfiuQhsIiSMywlj1c0/b
QYp8Ov/y9HUA5JEgGD7MFBx7ENEpAlgFGIRKDEsLqITPE7YCOHVCXsL5kcklX1w8P79vU+7T1mPA
irWDj9AGCYXoHbJnSXtyFmS+Hd1dtE1PZ3hDQztVDSGLfQqJDHXgaUS5qBVXNIG6EwCE7jOOUvta
LLH+7jOsZoJYQp07c95Ykx2sMg7TPsaBqRUlwhaeRE3VCaV0LcSjVsfnhCONs1QHaRi9CDRvfHHF
xeQ/2MLM0l8VBFMpesSduIA6B14GpRqfNQXvqQ5y5+BHLcRdBFkO2Yw1sIlqhRbkpXtRKvi/GsJh
AbjYeFJdsNAkAs6omecHm6s9Jy2K4H/ISi7E15+Jug9NOIi2G015/mLFMo+FqE2yMJplcXy/m2Qa
bEYiCzOposp24BXNBlFDtBLfqobeIi5zB7thXpNtDdxxOAfb00M57Z68vtdbwLso8arqNG8gNlrX
h+MCRzDX1AjyMZfiiqJBg/cbd9KSUM1g5KhezjQg2x8dalmv3o5i0EQSTc5vXSZ0pSpyFtM/YiR1
U2csoFDMysTmwKFEcwoWp1SZjn3jEP0VKYYHoMeIeMURQUGZKpty5facIhg0/p92x8CHyAYFbo3C
9vmYP4E5yy5tzYCgrUJ6VPD8AfLB8bOYqxJ3/S1h8u7dvnwLYiEF0mI+eh6elKZphQLznXm062Z2
Aq+aiWSuK9MYBP53u3mUp7Yd3w/6c6zwlL2lo/Ie+6Yl5msmh+ycuZe2BaqbXOnz9re8+raATJG6
OXhbWWD+V3fpqJ6UWSrAIE7N4dRGM4rAhAepulQRIjJgRR7gJmo8bPaWTYHu2zJPH5F8LeG2GqQQ
gtbITfNdLeC7bk/iU3WnbisYDybaxmjD1dpVteUeHdIbWEhxYZh3Wqa0Sc1mGWWWmZ0kIuYSqWe2
p11rC59ncBO3CC4AF/gob7HnWDUkMLLTNNQeXeVr1Qjd74yWMO1q/GmHEPdaDpkVSOqgj8aCf91B
Ia6j+pR4XxpyLs1pj6G4DxeZ5JxotE8pBH4BYg6Zj84/KvNRFu3WeAY3h55x387X7fYGsn4zjH+m
nFuxIQ0fMOux5cvyHwfdlHutdv5BRpy4zGMaPO5rvvVt0lzYfiu82554I2LU+NwXLgx9UU1aNQkV
XrD7ko/oY9vwUt+vJCG4go79pxmL7jQTQXhoNLlEpzMcSj3/S/VPwHCVRuuCh0qep6Yn+MSAt/dp
yZPA604UBsf8Yqm78M5pZ2EbdXULiMKGDm1NrYuOi33lrfjAT44Fj99umXBizhfL9vHo6xyqe41d
KMuQFSxLQEQZrzjF5/5liHkuqmxEY2IXlEOkA38MG+LMDxl+FPWqTPDC7lAu1Orz+LGQDr72wLjY
qYeX1qJwFJv7yw/yTThgo/S4Iu92gA2iiQcR9jfQTT58VaWchlwadU2jmpV3GlVng2t4/MUxFc4v
sUaUk3UvmoOeIvNrfc5WL/oTsvFNMmneyvquumgLv015R/SUGQDcgeuLFdjbajsJ9bP5A+ZEob/r
i0I+1uRK1cI0+yd4AkdFsGQ7yiX5qgqlkqJlCHXahTxD7bKt+IMNmUpuBfBuhJEjD72ND4OiFAvU
MrIAgLKlDDptfZ3tLAlu4h/UP8J2qH8j7/bZRUMt41IKlu2qGbwy28qVG7zdJC/8UIQYmOBkQBOD
0bHdRHd1T9gXhgwQszlCwUGN2jkpgLehgc6/+OFoBtw04pD/11kOZhiO30EtpxAI4siRoreGlUjl
5qKlpBdYG7lRqau7Eh6uzluSc0KLZ+CcSKBCSXqE4qmnBPNrNY7g6PpE9EHRF7lJo25KI+ov9AHO
nUM2Um56NomCSpkJHM2YHVZ1PsX62Omaa3sAtxrYrgp3XvZQoLTJX+QrUkhQCoApvYD6Wz02NBJn
6ejnqRviu4aKJxmLll0W/tqVvC/e1NZxOvefq+cbB8JEFC5eOwVGKK105oE+9gqJT1AJB684AGk3
679nCX00I4rY0d9C6O48X22jnOHvW6mHGIJDfQZu+VzKkmC7ljKKcvxra5kV2dXp/lmms3xest7h
8gA0Ctj9q5XDmPQQc7DKQXXEQp4qjM5k6tZk+d8lYwJq23rObudLjgRXx2yIMk94LWqvY6OUMFFP
YHXF+933Q27KxCEYXIjtnBZO09BKG4/Cc/Qji4unKjSmy0O436QCqOS5KmUs2QWsAXE5FP37JHX0
oUwI08MY3523v9z3I4UMbrqUmswnV4VjJgjcaJVhCrvaHxyY1nfu6YhPjNgiOrAg27eW9naztI8e
6F/eTVva8C+Qscc3eyOWue6+oMRjRnsBlvERjWhovffIvevdDIpaIPZUHEd1VWQWdB6H2d+noBJ5
VgQOEiI/ol8x59sWhchhMygWULTr7wQsliOnNrq6ugV0t1oiHrrc5T9mZx1P+/QCHM+TFml1vVIt
XAl+lkHftq3DAk9MzyUXb6T1QBUlQaai2J1f6BOlFWrSwYwXGjpmELIfSuiY7+NSAXD2YoCr1Q+R
ZtiZ1hCNp0ywTaplX2bnG0Wnke5R6E4ZEZK2+7vC9eyh+TvpZFG6OkNmU20cwp6uT2EtlC12bXD0
KbIj4Q4jgVI++fcTCI7iSlU6y876+5ozEA0k1oqv2WQ262qlfoG7opwXeUW+MepK3tCpNv2EZnwO
AlHF2w/hS3C0A2NaqicPNRMR1lEM2rSoxiw6nKHdzo2tqyf5dVIR/amXJkmZwytFAcFlNq3owPUX
9L2uqiOEVEWdZgw2Q5XscJngBCUb8A7xvhy76umGPGtULAv8iXeh7XHk1qO9Wob51qpRK5rPMgVg
AA5wdVnfgidMDg/gVN2cvN9v4zrlqa50VcZv2Bb/Tl8QGASBk26cCdqvLitAY2cL7i2a527VhvIy
ar/ZnYRFnYsgUV3yQuMKYD4qJRRY7FNXYwkMQERfY/Ppp+/5EK5k+lV9LlLe6yPP4L7whJLhpL3B
fQZl0jsS5JSkUSKV/pJxrsvqSXr/EXwW4aewxPd/kb+4CSTD3Dj1rTguWyMXRX93+4RniTAAgViy
q8Lwj90vkrdYpxia5uf+2XyZVn00GTYqH1uISs2LcpWyejUR0RHwPFHxeEuuQ6rpB8ImMCS+YH20
uhxrrgBRZVjnm2FGC+t05Zd7o6eOF27vfs8Lp/5hgI8ZsIx+M0rfYo3muBhxe2g1L6kAPtjs0LpB
S1ht4VSEd0FHAUHj2Ri60okV7xEtcCO+Dn02CCHXIHoWe9LdiTOuF8E+nQ5jFPcoarCTgmGVd2Nx
vvCgGki2Sw9P9RRn0zcS0kWW13XrFhZJiyP5eE9otBr3U28rUkxNF7YdHi/gbVoMvOyDVkudjcwh
P5RAc5PcNa/VoHqFobPbhx2d8kyOUCXNut908rQgfxXMfE+AkGwdJgUTOdZfrWolIaN5wy+F3iN8
bphWbNEoaa3FK34mvxCAtKyjGRT2wGmjstZ3lCDROeFZ5Gk/6WvDvHfUxs3jvbnN0rFFbprxQBTI
AfqMndfALflLWDV5+0n0Kv4pzmsto7XaFl6zQuXCCoOJClhf4aQ9SmzD0s5eNzd1pA5PRa3vWSzj
BFw7bRDo2q+/qXQMiH85A7yNRO2ghr6VALYXjBAwZrAgs/JWePJMT+OsKJ9moU1/qPMuONhvRK/n
rrPCTDOEwZHl5lVIU0CIZSOxQiY5haRkwpWo4WlXqGBvtD6kif2TsLxFb2Uw01yNNWPYCeesVsWL
ExV7ONAin22SAxruMUK0BrvkbWlPv+irDNEaDTKEJChdCRG0aEpOolwB8DWpnC2DPEZCE+elJ6pW
i4vFyMca8wt8xnX+/QZOSQG2lXLU3Y2lvsjApn3edBta6MdjrC4Wjm9w/Hfo5Qr5AXJZ72icijaM
WHZEy8Wt6RHq7FjYj8IUiKWjAonOvWRybI7GSBUTD2bkyHbMC+XoevxXwzOS3aQ1BOtcq68VNTzJ
t6EIcB2m5WLZ36KNHnFQW5+uU90MNatioDcLYD1zGVEqOoUTRS9zQBcjZvz1D9EdhxNNbhDNnzqq
jobtkprzdaaxTzVpdkug/gRa6uQCKMNV7clLaK+Lc/99LF7R1KbzwbuRYKG6aaZWGPaoHcm3rPUX
6hQ4OvPHnPwW+zvEOup4xmoNw5qCSbljWGmEpRo7WPRGFvT/y2GDaXuhAnWAoH+VGXhSSdRZrr+3
/FIfK/pm1mDCNiizgI+G1IuYBGzcbzZv2jv0wfe3GL3wzFbGIpgcQnsKgxM9KliJZe7ddNO0a/nk
4vIcI+nJQTZUf84moT2H5MRNhLmIRArN1bFmgm51Z582sYn9sqDN2WtRnb4PNGu01Nk77oCDu1Mp
8acHo0n76FR9S/2TXK1fK8QUsj3exYuto9LR7TK2v5DPI4e61badNLtiR9tG296aG1nBktUZZSfR
OjV6WHoNOKHxfmzrWFIXTWEOZDJm6tEjoGQ0DRY2PZyjtUzbieDx//ko7UxQeGKPUMrt6v3lOVw1
mLORi0VCCAJN8W+YbRc0c8nILbE0+aN4avIGQN0iftqe3JIr9Z+lf0ZqksVWMD6+e+fI+1isXnUZ
m7glcfMQA3touuJ4G9uNO9a02GTxdihWi4+bWbFBw9LDBP+C8fXE2znyF5eCvirajIR+Og/WfPkq
i3s6S3HecdzxqeeBg2GIXg7tpjtyTCc7gUmk/8CzOXa6I5PVwF4LaRLT00uTRtAFviH4wY+mxApf
yCB4m3x0nFVBJ14iMH2yhfNZ65f1/TIiUH8kXJd8p2FRRiD1XHr3mcU7xFMGemEuU0SPfKRuQDWM
dvXSnvpWBNmFNxcvYVJ4lnkzAwZUqTDIUpSEMTg1iGAlhtT5TPiGCRD4qat2Lmghf/hBxnAj/a+z
ShLKZJtLgsnoHtH+laqolF4mE/RXcMric5MjAwIeLFXUY9QzTtnB7Buw4urs5p9BES6qlT0PiiFq
DvluhjGz7MyqrYDSs+vjPyN6xhfsQ8KR85IWRAep0sD1bFqTWjucwyOu9hFhG0ONI4Lp53/RxzAx
S3uBvdO4euhKG7YLktZJ0zM78iuyu+pIV1CZqDDB3NYd3+oOv5xN29wXoQlyrALU6dKYWWJ1RLvO
VToNQufxqW+OABOxXib5wUl+1LGzyHYorQ8JdKauPEU4gHYjSTcrPegR3GyP/sC+yrjy35g5Jxtc
BXD9xwm3WxBYx+CKBKxClNmCPoU3fTl99CC45DSi0BYb4GpmJQC0uLvxef7EDbwAbwrKW1HtfKpA
nNhMyH6Jag/OqXuCw3YWERI+EHzqiLbgLBny8oL8NtiC6vd5gd3dyYgZGMLONVxk6r4Ni5yFwsiQ
9/wK1TW/P3W0uMtInwrtG2AaOL1amMGZN3n/HgLB0sh2s8GOKRZV54eaFhLvlqduSuHI0uAAUNDn
GpzUlMNHCyCEDPD5MJPXiG1NI534fycbSBSfdna7pGVuEb9Mi2Hoago7tcv7Jgpog2fQBk73gyBD
VmRENIZT1e2pblz+9AQMjqNtMR+wID6p+zbl94ASDGbN2cSMXkGt71T9lzJLp6uu3uABLqhgq8iv
ZHxgmSs1R0hmijDCFzx1CLCux6RUaw59HjbW6CiwaEufoj4z+P4hgonlsbc644lhvb3wV25iI3h+
CvuiRsDhfiilf1qW+iPtlBu9LUHV7qxl444oDZTLKJph6zQ/GFY8F3pC0Gp9EIV86eUdl64BnVmS
JbjbwX6H1DfQmFh2B9z1el6McAOkDPYKijQnOh6mj9BgOu7EASD3htcBNPw/jKc63sHRFvNeSTUt
52pP04TE+mi0Xg5gFndUzUr+/2GoQSZRFiDpm8UnV8FpcLdlUHjVh3x1s8D031lLeYs2skH1pKmm
IsHYNkeXrQs4JniqtciqBCVE1nJC5Q/FZnwYKJLQaYRIt0C9BdAptZ6/H/vFQqFvWKgDIgxhAiB9
EOLpFsxeX5t0+TPFGcg1VkRsnbXx9dnuyEii43CUY3PHHZq/dU1L+5ykDVgJxrpFHVIfkjCxk+sS
uw73/46gRmTDbt842Ok2R/dSca/ZqioF0tkKF0PUPirtDREVgeSuru1U/HdHe41sUdnr24cUZ2hm
0Ir/UYKESuK7VBZXWK/khqZjHkHIV4xFhBllNc5nDoklzGXoOzgzrL786eASyD0gUaXsbfMkcsRZ
85eWD4tACCJa7stHLKd29xH93SholHr6YnnuULoe2Cy4b8d2ghT3vHPpXW1CCMsLYnd5NxEQwWyW
1ZnwK+DHFEQHRHCKHHvFXOA/43lL9jtEkSaHqW++ZrNaD6RE0bufoEQ+cewAqnnfVPbyDFrkOaNE
lvR4vJEzt0ZejpG59T+flGxuuo9NMsYojEg220tOffItre9m5ENNRRdQlf8oOjtU+9iowVsDHSAp
NjTFNdsRXKiUHrdtFAKNp8z5s6BqT2D9gd4egKf87vi7fF5VIAn3MabwO5thg0dLl8b2mNO4CYcD
z5SCE5SOMMA6LNXG8PsMNS9+5ChOkl+GTM+8ee7rfPac5L0aWkdZQdSGlFUFOLrUYv2pk1fpqu3Z
7A3cXzzQ2ENuR+uAPiXEURirw42ymuXskA5moNJvStnE+one9IOcINPRU/FO2NXEl+Gd84iV0+kM
A0VrMukJQ1yb8QFPgseMPqgg+DoI0S9/ODl9QdiQhxaj+uFh3PXOXTO3b5fYimUO3SKSBc54c6Mb
af3S23Nhti6i1GwQhl2DTu+viUmMafC4zA9/AAPL0RSKN3krLE8ncvCM7UyVks8gvE4Fuz+HedwF
LPJ+IKjdLtRh5ZT3+mzocoDkMhrqJZg4sseVTuoKiVccaVSki6nQPUbGdCh1GvBOxch7oGQHK1mO
iLnN6SjO7YDWoCQAs2zIbmJ2yP8PvRHWzUHUthfrKCmIUvkx54ha6RcChLgFyVN0FDrmUmbmcriv
o7lNjDWXUuC9op28BR2J8zQ25dw0S2Cke9n3tZ0xfunMeB4jMAFwqUdjeMsqhWIrFPSh0644XNJ7
Un7pjfsJRzUBXpwAQ54ki6kBBSPnv8m32cqCQ5+qRYKfXLGb2QbBwN8wWzalxT2aX4Mez5Y4M7MW
iaMEuAUpb6mkyHcW4VaS+SIsSRmSo1czE5SrTqBsCMDLhEhSPf4A3Z2hRNeV6vhl3Z5ta7etlEVw
ZOE3ti8kcbLUNkoOyZd65nRPX3zEweeot+qkbY/SoXCfgyMfe7SY5xAWjfk5oqqSZ+ej+3zFWgYE
yvQNvvQspQJuQcpNBhD1W1UyauZbf7ujfbOh/+C/gl+FViUO3j6143HMORrQ4FPADcj0MmmJc8Zx
KuNfzoMRwFG1BUj9ckRMxEqJ/uVu3uEFxBm9KEYpOj+pk6MvuwzBvjEydmrEWM1Eqj5ajDTmR6vu
7vqTewyAWmpZU013pUPOYv30MJPU9P0Fmkon162Isis51OY7cNtihKQyTG25oOUrI7/5NCtZDbyA
AW0P+YTScGKL457k1oZcyoR8ZwxnuBVSHLSYKvlVWV9ckZAlDSq2omwqQC3wQIHoMytStbUYJJD0
0jfC4W4FupI1Onpo3l3BPvSTiUZVgV7fDaHZEJNm8FAIFBY2SV7AWQ1loxELXmfz4jGLdYjNReGS
q3gawWY3YjXVryV3QT0StbkR3ArJAPlOT5hu6YCnh1jwApjwMCfKJFwj2pqzCWpUOzhMrKfmgdM5
Pni11hp1sylTXvgfpA89bh+AJnE3cubaKYU3Aad93SGlKxWpnsSlfQtwIBarHffK1A0XJLJ/kDCz
or5ZJgjRbzwJ5ogLIpHbUdnR0PNJh+oh68gjGajcxDYqn2M6pb27je1SqytfEBeLVnHo+CeR4LuG
lOMbP17MjZmY1p/8Gl0P0m7WFCwTkNN25mpNSwHpf5nWbk3U0GeykxzHRy7LOocXlzRfNv+USyiq
4abLMaTShSAHYEL0n6cEI7dYBIc+uxP+AbOl9BTmqbFkE3nuflAQ6yxkpTAav0l+hO1Pyeum5Hp5
AGGrauO6j6jHrTD1kYIE007hcwvaptGfyjvohpsm5Z/4UpvL8+oTtRxXugI9vsj6LjePe+78QFzf
VmT7zjnIsZMiq8N5zMvqNJvzKVTMcUyXvuy+JansSKSgby1W8WW/W5KnLlS1jWPBnx8E9NXE7UFQ
O78gdUS+H1FXGqpQq4YVzlL5WZCRB/6a1cZ6/N3ir0WW+Hq65BTv0tI6v7JWawTfBXr+T4njrRpR
cC1id+5/TK8iW32rlGhgYsFpqwfTn1Jg0Ta9nYYug0AfMILzz4kpRK3REBGd36e5r5p0UqBTbyr4
wN9gVb6ym8fWDjo92VVvXS8C22e/Ns3hJlQyzxyQbcltglYcKt4GKvrmBCjRinq0kal0i+4/YHT6
Ct3Gl9r+0LyTvJ/Ls+6s9Lh7G+QOdavR1GaJuQnbd4i5BGLBQ16EMDSCXYIipz6yOuS4TI+/TGQe
+L+5tBNhc0K/Frt88xMuJ57aM6izAbNwKu2VABkI2tHVlgErdIHVVFuSkku5TDa0PsOf7gtQnHYf
9lHY8MJ3RPtiLhpuLxBrsQ+qxa2CcOjIAivOhcMXzTYaLoJpQPGfSVmJ0uDqXYDfOCWkqkbnqydz
ITSzbF/rw0xmwAtyfh5Zu89n4NJ0XyM21ByruxFEO3qQqL0EclgFL0zBaZIpC90klkvPZsiOQO1v
KGKAK83dZtFF+HYA6BvSfJ1AyrhQ8ZhDEfIcAof1/W5pb0BDcKDb6dfVKE2zpo0SM/AP7BSlh4RS
Vgvd9jS4SEu4irRZZHjv7bmBMzw67T7CByhmEuTxuIROoRiJkKp7xpEMT/rzpG3hlf4r3z4yBWG0
/qrt3LroYrTHuv6tzMImf1KyKuLGvUfp28Vc5EWiHL8X5/co8aRqIDIUTukyvzRfIpyiqCOZIfUI
VJC1IdSim7l31J/ZGAEXeZkcXwUzwGW7L/BNgOVE1gF01KusOA3gdLH9wFIxE4QVYsr79mLcFAKR
Y9o2VMWdmssDQOkNoXnv0LwJkRUHQXCS8atIvpj8DuBF/tXqPL8nDtqAxFRN16g76nPXb+P8+lDI
1vJ8jh9RwPAXi8F+LQfkc5FRHg3xCPGtgcJ6E4f4UxGB014gcXLHcsVDo1Jwphg3Mdd+Eh9rwka9
ka/1soFaUPLNE/L82HxjgISEoDd0LDk6fBsxkodJZaO3LuUgrqyk45tR2GG6RARYRqv+5nUn5LvK
ZWSWDErd0B2WoNUsHK8WVb6Q9QOYuoc4RxOfEdZ1FBgzBs9zexzj86INL6MmqKCy/v9Z4ns9CMYZ
SwIjUC4dZrZ5OiUeARGuLLIz51ICRvx2vD/N2UuA6CpAHSnlMzMnLXf0YP1RljHrxgnFTyLG6lfu
gVO8aWRs/u98BC/mX/QtaU+LM5fPQgmfutvD9cHDux+6YYPqx9aP42Ad2BN0uuDLwYZ+mSE/vomc
D/bdLvAkEMcfrPjDtev+kmjJyVDer2EsA53be7+MOmgtJiCnEizMfphDw/tSAbFtgWwYWay65l08
W/I3Vq8poghpp5yvL921H8LnzGioFhwZv3zLl2K6IvJAGaTcgy1khGH70kbQt/eL69FIsWNymYNd
8QndqdFTuUZJIFavEL5yrrSubGGz5tZId3foMIaugkiI5sQeXergOt7tNqYBWPjfrMqNJ4ruRmOC
95eOyHJOnDsDJ0UYSwU64BaZJ+GtJZBy82C1GDUdWtgiFzRbdx07WdFCU9HBn2dl3mPCAvHbJ9iu
NszqAi/Ty3RIuE6yd6IulYom17V/59/q8YMZoSerDHSeTPh+fskgKmn7lnI6i33cp4VGw4SXLVro
fKgAOWdwfwn4/0Wh1ZfItYIZMtAQC3TViTCdez1npxYTT5NFkQ6Jda7uzffxtbI3nOZ5RRz+MoII
D3XQzqgVoHyOmTRLJyCjOFfI4vsw23LbK72sJStu4YIMA8lqrqaeftxLLVPSeqgnTo1Ntx7dYjZB
evLg8l8PcZARy0hI90Vhagsr88U9C0FeNLHDALfbWfRYCFFTkwsXoBy9v3NK9UMxDe8OgRhx1OBg
CNmcvUutkB7EgZBjboJYQs1x/3zTfHk31JqmEq7EuTD8Lb90eqEN7bYhKgG8gZeo5NSV1ui57S02
sKQqaHdLKEGfAOMgvec+EU6Ad2gq5B94W3O/P6DSydjgNLwUN9qgp1zI6qXahMpA97ekQlC8Jr5U
H6pViYERSlxwndwcs8HJI8LkRp+2foNFLlca0qv9bNVuXZL3M0Z9N+ad54wzSq72W3yrky0s2T5c
5HdpyQcthpdCbHsThWDUyrMFQdui5DeajWH9BS8UdToD/QvCU2GDlO3WVjNeTYCn0NOVG+0UWTXo
y+0wNp2Bzc9P78TlyKlcmuFiXtJzbE0I5vUNEkqh3s3xwMMBkkgU00OzuJpxPOENu0p7r2v3ZaQb
Y0E3cmvBQ8acfgkSHK6iKFmaellBMvYQBazOykpRUfkAZyS0y9obAkgoIOT75nbFK/DDeL9+WVuN
4Sp+U5W9wZHANOGmv9m1y+EEIOdO8GCl6OZbSWolaTddCiOqNhyaf/zzgwS+3vdkwNL6GUwNzrDR
yssGbEID6ThKBaCks2V1shAP0kO75I07ljzG5nt3IiiiSjpJWa856J+UWhKVW5wZN1Ezc2ym6mTI
BatlST95hkg7skmJupyWXyC8HxdSA9z9aAHOLibXQtW+Yc60HQqA3aRU+P+jstbFJ/vyxO1hs4gO
Z3hN7SOKt1jZHkzPxlp/v+Yg+/0tRoDUUU/d7kfGpu6g4sR2KRbPUrsdd8JY2oxUgO3ip3/7Mqry
CdxcumKsHhgTCLj8DYCY7/WgvKzjxRAU/b3aWwfKFT6/fUGMBpP57I5GB+bbM0Txf0deIX8VgyWI
Ck7cYMHGQjKQvFSA1VwDcq+o80QtVO8ycTq44hOWac3Axp3eblZki3fhYi9hOI1aUlvWUxVgKfh3
sEsmh+6tLlTXMth+ABy0739zVp9tdJ4IDfbPMkI4qtLhd07I0TpI8ne5FAc1Bzy0jmdXxzTfcAuJ
0P2sMHiviQWzr9TPq3l5XOClqbaIra3n5AYUZWpWjT4iLZSU36SZhIQuhy1yrUsq4p716HqY1BMT
6K1+HzfXOYL/J6ES9D7Fjg33LZxr2H7INejzxkSb7XipS9BAqmdfob+VUYzcmY7smANhnpXzQYri
x9y+GZDSm4SynRuumVGIcXTbRWc/zhgGKImQhZ8MXNWDbbDBlX7foIKlE7CWdX203PGElCr/QR1Z
g1HOuHtSHVuxwPZZaeaQu5w0QBilNnowFKmo91McCJW5dNMGo2ytGDoi7KFOFR0pTJUPBMbcQOI7
2MSatZs47uWg0lhngKhmGxR01J4UbgN03ABTeuakdnyxpLecQLMCgzHm5+6R1Kr5Zi6OGcAefAb3
dUqk5wa5EI6CePEf9Disb2A8zWQxTTZ9t9Iy3+McpxxdJhVXFpjuElUa3mP600vJobu0e3lKZbtu
T7lUk4pB/YLd/kRALpIZV/UfuWNSnxTJqGNLn8AmqUWy+2tet3DT7P346uM+QFtytg7prHTbVDmr
tinkhMW5zJmjvsJdT6LIavYmZFLo3YtbmVybI8gjH7+vLup22OHOJRcFUWIbRZHxh8AMULUo1YOA
6NDhV5R1+GCZB0l/1KEjGKe7KczCYSH6B47+n20APcnj5tDXkherXO5y4eI/XOe1UiC9ee/5Je2Z
jH2gXWGbjzHsqXaCyViYGjrQ/41gipOXpPfXkam6vjBBcWVgzQiXhiqvvFbnV7ujSBVtGqMiU6h7
MMJ6JnYHYmruW4xIx7MoHFy5LD8Ni8UIcungNw8jjSEGQASfy8R7b4QV8sgqpMFCOm0JGnsalLUh
q3yalaGmmVdZ7UtRZ1vdyEGskLKD3xioBw4bKzwJpAtmpgPL9Fcl220A7kb3PWXe/fliae86Zu6X
knDws4URjljwVBirrL35KHBaa/VCc8eslI0qhwd4zwbOTTGXAff8cS//mUIdJX2Rxk7i/JjiALOZ
CForhRD4i7wOtgxW7zROVgnC4nmAqWuDku8KNnpb9aiA6jBxujv+aUYX1OKEvjV9B7QPvlXf33N/
LnlpwursMB5ftZ2ECQZvXzyEqHn9V1I/UOD5BjhERD5m4Q3V0kx3EnK50NmNQ7cOGrg8Co8bAq7H
kilUl3j0fNUYd0KaamPZLuFRXedkqEAaCxLPHZgvQzeaQfq15oGSu0j8yio2WkmmapGoqK64dxGT
RgbIVe60mOBHpYaVN0ac1oGrIhmdWV1dlfo1q5ZOohHADxnDZZAti+Iu+jISNSntC4nfHzUX6m7I
x00RHK+Lbl0CDFyyHMRvF9Z6UfAaG9vmF+Dng7v6P1KhZgztRterENyYCQXM8UFHuOt5S8Jhn/Vi
BJ9SkirBbvv9uz8MQKLSdRHDr9KEWJ35dAwlCXWaY8mdnBNjyq8vHArQpgiAmQlAjwkAERRVWYwt
3oER+KZw+t3GQGRkXdb6nY/8BcroczsicCmT1vygVtQoNoabGuPwHsA9195eCNjxJkpERudo89uo
WLTw9MMeaZ6bH5oD8s4nnhhFC6V9I+SIOyNzYt5apY5bwzx0DH8t7p8U+4a4btyKaI2YLbJxw3eI
2jKQKY//nTEDHbFbVJG/ynAwLnLVzqyRrqOIW796NIAPsX0dgJjhU7B4exRh4k+bf5B8TY0RTvNV
T5CoJmlqRYQRmhZe3rsnyPPXeAtiGiTclZDDt/G9VefFBlLhGHB1EFx+qIOBEtwanTam3q3P+WgN
8J9rViWp1qQy2tOoqmlBVDY1P7n+Pr+VPCoeIMsTm6Ex0W9zOgcrLqoTH1zSjt6C1fuL4MEpFXZE
nq4AvtZGpZjQ5h141zE6QnA74J5Gr1BtfZobrUlquB25paqzuR3EcotPHn6GvEaROcjrEkiQe1pY
MOWr5PBcrXiL7aYNRt3Duuf0yvM3RoNDmmIczHedbzycQhoH0pej04IslmzS8uWXyjEIqkZJLx5w
KRF964YQaBobiBngN7MK24ufFWpwn39mMxkL4TaFWlubPG7QUECyXjTXg5xvIPENEk0vGgE7TwyM
CQTGFY/ZAd4ohBW3qKuRddNmGWXxIyGwWKhOrhDNGv04wy4CSfwuRk5P18qB3zQC9PwSRkQnozGb
V449/e7VhwBaTAcTWo0bEyYK8Fco5VgbAogMIoDmpqw8y+zmzk2G4Sf5Ki/8EGrpUGaa+EF7AqMY
rl27FKK5OqAMf2MVewFkgSQKoYXHpMWpO7IkA7pbn2Ho+SZPwK3GXjU5nW0GnNlhk/EdjClSaNs6
3zuYI6SE2S51P+N3AQcbxgcgZer5V1g0mrd5qQFVV0Oea/hU+UdaTuDXXAAr/JZrbaC9QLbkm8Af
IYXAZUuA0qyc2RX3paW2lhAHnfR/pwuq1FufSDkrZgW/UUbojB4PMoksKEWvB7D5Mh6GXCmkIcy6
goL4cspk/0ZdaIdprs5LZa/WVfYIGwpjuUJuOk767wfRr+lDllKbXm/ndpwNdlsvAR2SfnAuOkj8
CYDCQxBbPZfaf2Ghu94NegL+/RYb93hwJVY71qDZ3J8nxAYhvMrbbQNOu3IW7TCLsUV7qkoLgcmR
iwTpo/1yQKEh1ViOxxqPJdkRudFt1IJod4ZEdI6Nof4rN5+7cpireKr+9QpRPgYMmbCzIKKsv0b3
SbPC4pgNTHz+NFHwzbHk7LsMUMuQJYDMBgXcwUp5jXCodUC3kREgABzbERAU1s9xGZluIxc/L200
JXwinaPtqKgvLF9hvuazEzdIKNlozCdv4nf7hz0aTWB6zciTWsv1SC5pvN9drME2pWVefcrkjRDe
VKjg+d5hLTmHPdvV4yeG7jQ+wosl04iYXgPKnf/9dcsde4e3aJPlBmhwiWdhCgoMfIGb7e1pcrzD
KGFlWweIQ3eC1IxjN0ruGAy4L7AANMk8Zkx7fDhNJapYE/cGtutuZ7tPHDB1Bz/pohhwuH3cey5T
SYqMkSAb2HYXXOW9+/ipMgetUIzYXirbamXRh/LWRWxu6MGm3AZZL3gv8swr4Ku5C2PLKKy2AuKx
+0tr/HF4zkQbX6suZto9GNrqlcGMW2r14Vnp9Fhb5CW8RQrcqDMx01R5buBT2Lvmb8hzXq/6mSJP
B4JxpUVux1i9a+l9I937qw3WUR/Nu6Ix71zAtVMMZkqDniBNCWzJwiLnVFmacOPHu0azdJBjmFpb
sVMb80cGR4gPvtJIv8TkFuLd0MDiugLGpICTKLiSKEp/lZer2ea9jUaMtEE655ObV2rE8d/pbhM+
+jw4buFc97WsBMRKXk3SZGfavrIuDDHXsfrNVXaIuXQlAxHOyy/WJxgRQ1r8Kre9KYwJU7horIum
DQXTcTa2LXpX1/MqFzWd48mbDiF+dpv5hY4mInAMxJEiWkMV7SAXszJhaxVV/5FTJoRJdqnhKFuY
VBh4GzwkejfKpZCvQ2zTsumm77turXgf4AIV+DDArOVXnyGtGet+7CTv5U6OIfYWHYxBu/dZcFvm
FbemAB4MdWtkso8dxdn6YIH7D9zPnLez2l9wsljrSp4yMk5qdcwiz2r6PMVss8N7dUKoVvNEt6QM
jaxULEUmELR7nrnVCsh8DxQe+eZ8o5BbE6xM6x6ogyKcKvN9pPvoG7CNTmCPrKhHrcfgOrGIFclW
Zw11zy6xgSeFKILIxIflMkeDczDyitM+I2YWoq6B60XSu8uTmbrie6QcobHwkHfupm1gY34YJNxS
eOWTMuIJw2e7mmtgMMcnhsMrLuiYhFclB7goTQyX0SIADgF7lD2YmYXqy85TPHoIdgNrB1mIFAK0
KNtfmcKRMr6Q3W9rnbOO+7sJ45BJbENuvautZgO4Zdo//ehxi+hsBGC1u9JUhLdnNGMQ6sSPSLPE
0YhhS9+R3+kXWwgt1PcP9miIQo9WDe6vTaDaVn5x5y2iq4bHwlOTYpK6wue6oe8gB3UA26lDd6iU
bNQS8JtEacB0Z/1kBUGvNBlBypmMHGgMhwLpLfMfSPzWHzGL6feMiKXcbtBAh4AQBl8vh9yrr1VD
Gy9nT6jzjeKa+KGN0SRzSQPeEeHWkkWG8smy3Ycncitu4lccqP1JHRxVjmDBBF+EYdZlFVrHgKXi
D5IyaFyo050ssHTBCnFWMKKCmncO6FvI1G1lG6U6vyWNPDUE8IprYauKamFbWy846WZf7NkQtLB1
UjVAF4k3QndHEx3E+TGugWfWgmRHypdZgHVd5ODXcE/69eUYkK9Qvnvabhy8imehCl0OGtod6zyG
L92g1pjEFS6Rq1ZUNeHt9skIcfY5xt1/CrbcEsizBspOroerbhqpEejqwWlYx3wDZBUo+CRmUsnP
NTQimqTphpqlOtamYu3EXq4Th/MJub873lDeY3dvS0w2kounA5VAzxTKfdYEEf/uJzV8r9RXm3UX
RJOuue2E6qHtlE5MpWCtByckV5ZHiHkXxoreVyX3SUK/jJETyuYHVMvrWhe87jUkYI98MhfumBiD
Qs7mLT1j0PCpCqVLg44SwSpx86sW047qNYIfFPj1RTspC/+oy/oCE+Mgo2tHFsTbdzYjsgMPXBzw
Xc8L6uy8ml2FWvsCG2Y8EsmNRdG1yO6KURbrygLC9CnL9epJtQevzyCUsoe+cdMRQycMIj8pG25P
TCB45EbWxaTBgTpWvCKr24GBaavJSJkz7/BP9bDx8ZrZkG6VBcZrWvpHN8x3+MKWb/houkUIZX38
YTlyb2oUa7PYp3i3JeenGKKm1YTLnAK/CmdID8uF7sT3JnVlahXWBY8Z6YQJYmAezqc7z0x+uNeL
JXR+6a5nVFM5Y4NzryweImip9yz0KcEcmZHjvP/JyJPIWe4CpDxgWwHOqbipzh14uEo5LVqpnTMN
XVIRe2A6jazRHRDzhaiZpD1Dq8isGsV5xxFEKsk8TK3guoPDwAbdm7vqcHNWcF/RT7OHMefvd8TY
7HSylDjR5XMcB4KVnv3R7jHhtGxvVDPoy0PZ6vlI3hw2l9xVGsR42Kn49h4JXKMQQVFm8Be2EbTX
hF4azU7Rp4cgutKp6loF8YYG0bDEycd49fHs6oaRdz6ytI6VmyStdgmxmM+QMDAjYu/MHHK3UcfM
cejG8IqllswjemRVn8iwhXJvzfW6WhkXzdIAzf07d0MD80jzQSO11etl0Uyo5KL38qi1jMmFwRF9
gkPgC5ETiyHP4CbUoZx6GqvOUnuv2F+Kvez2AKO4iZGlnxtW7v2uQzK2KvQt1Lwjw2CLcrIAl2on
DYhyP38KBB+IOEpngFb0t9Pn+iYtMfuVQK34ZgMIfvdK6sdHq7B+Cd/Sse3guogoxwqLoHx8Ms/S
6LNt/ej983oPTHdqJTvnGrjOdl5zJP/xyDkPpiTMsaGWn9wY3m0mWGUPU0wbk//P0F8SBrrchsvc
V0iaASwhZGJGFd5YzFrOvFkL/idQlyuUCRiJQfavNfTc9Qmu8kPUBL/Oxf1cm2vBXeZ9zjbJEuiM
Rw1VhvmFYvY53r8qVsDfwDHkQ7qYxeOUaZgHrM8SMpzi4GDZcLUHAOtwQO9h6PZcktiLyxYz+8wm
tQuiu8xDrIZWPUjwUo0fRB8wcB7smIwY7dSQ6dBITAUuxoqOwnI8MghCVc8sdbTmpRIPx58aU0jq
4u+DgpGlGtF+CaDz/IwMCAk6wNl3ohN6NhdOW3iCBZts9UDUD/HqsoCcgqyOua0qdihxvvxRRtEU
miDVLEVHIAdvBkKN2+DZSdF3tD4ox5kXE5FIehAK/c+Lj2KBWQXpv8V3rBqsf3tqw+0V5H4zQa1Z
Jq7/JmKTSPrSNF+2AD2R/LrgxP7e/SGOaS/ZBxkuMUcvn30n2g+nBJn133LrwShEqVLf9K5Lq+ff
6f7nGRAGb6PjCg/5t98w8EwzXPvWLiXxUDVBlJtGv17RWZeSk+o0gwTk5c7wOLU/+fSSe9G4TThU
cYDRdyX4MtHdlVnfxlh+azSWAT764ddqQgoFMViQXQWkXVyQLWGKd5/x9nkpmy2OziYWn+snUitz
+7r9OumBeD106DA8eu/fs8hTrmY8GJY7TtXKpSNpd07mOnqgiZl2iAKnX/gPY/iugQBSs5sD3L5f
Zj7jgC7/5iH6VPfubtEgEka6/LClbpSA+aVGDgK49PJEafVyjjbpElqDVSTqNR4weKrd2r3qx55F
wlIt2kQz8whjAAbbCV6EJBM1E5/pSI8pmKXq830GL0gY0+2yaDzgLtKUBKgngmolSOYW1rAIiSnL
h9K0OpTh/HZCoaqn+9zJIfxsP7YbmxSFmOD8k6T08JhnzGQeFkIUADKpzm5zJKEwacZXfNf4GbKP
cx4ZMa5kosvavI19zJQiCnjqh5TqBy4tt3fPFThxnf4Diq/sxCmWU8fiiAclR+D+dQXHNxTGXaOm
OfAbUDDvJLdOg0B6NPMHfklCDfJ1J9AR86r79CiHAO26U4k19dqL0FDecLoj6f6B9JTCxlVjlVFD
LNwNsd7fKYcuIDNBlq1p+KZ74COPpMRPkqalYd38TRSla7u62Krf/RKdEu01UoV0orjm5Pn9ogUx
7h1ZC65tJnI7Hb/JLxcAaWsB2Ln8vyXKNKhHZF21qKG+HkOpzHC1RV6m6DSsVYMerrkBYW1MzNbW
NO/kfRHNAr3DCqj0wgibZrwZaFflBlXoQvyIR0glv66/zMy0KSKDbc3YfxPwLZQ8zmCIpLDyII9I
mYPGY9StD4suOsbe7U1MgDR/aLJp79iebSiChEtApX7cFVFsGMMbb6T9ZIvQml8L8guGF1bNnYgb
W5HX9bqYc0lyhIVruz2BWlzNwLkRYt9o/mbuVdFQpaA1oygPYt6H9R2zcRRpOuH1SAgIjr+vJVxI
DDgDCmhZGArCzMHjhR7jI1MP23dvIGi/qqWRO1BDKfOldvyguFTnIPzenbYpMLaAD8nWh+kjyy3R
SbuLB1NlNbMpnKBYjfgJZnmYR+QEUpvbWoeb6vXIwwDj0HaCHknFIj/kfl3WWdc/h/GPVnhYihyz
0/Zm6zSMTRREDjj95pVWalDBJ3H1fqNw+HyrHLwcAa0osE/YyNEKIdzmMHO9LwDU2xD8e9OqKAvv
u0qoT+0eRAnYt0n3k4Bnn4dvkS9JAWCbnEVLpCdIRq8jltMocZPJDaxAs1ehwMDSRSANlvxelDHT
ra1P0fxqkVMA5Hpx0/sTELu2ArpzflzDiJM0QNEb1OT0KiSmyLaHBL/wJ/se15kLvDVzzFH1T2tZ
7NUCFfG6Jb129tzBUTwBj/3R8r/N/XDDYPHdYA3X2kAOpe0CYpRRKpWyVtgsz5hshrG037E3kZY3
JcQKhSOJDJy6VxKDYCDm9Zd8HRpFWHW7L61vUrDkBSeh5V4M7PI2li6fKdhcsTrHGOeD9CCy3iVa
JIVITkNuF1L2CXOLBCziLiqH4e79vrcRtUZHt/BAXmNEN+ve75zz5M+9Y1ufRKIgXRv7roHq3pBk
QiLq3ZzgwBv/F4DA0vM8qNZmZKh0uJWrUaX1BbUQZJtjeo6nOYgwwm5Rk8IlB2FUs75D4e1gNbCR
MmHP05NgDiQZLOQbGs5c89bjX+c7sbPOe8NV+IVjD3SuLO/F/7i5YwuwAxZfTtPNBw/MIpamYVNV
zvmP3oD2i483qJ0LMoVoQ4bck715nMp6oj3D+8DQvz6ZA3dv3pRCBDvSVF0CeV72DybcBLKAk/e5
atevBH/aLWzcaqURGTb+UJmm/PdRILhm1s3ZjOkKb5NG2NC0pdqh/Pb/DHc3BRy4yRdCtdZPTnxl
gHlLYxpjC4QBl2HhTZtqfU9LcXqWy3YaLbh8Ei/qRgINZoDJyhEV52Oo68ijUxK7OxTw6P2GVFh/
XLISubgEnU/wrxYES0K6XmeO22Bkma275E2mY/qpJx/kkN5UA+qGAFV03g63K0CZKt4WvJjUDTh9
V95E9WBASrd47glnVhK9DNKwOW0aQfGOKdTvd5yb7o6b3MAqCHB8jn5g4qT15BhWY+90XNmCU9Ex
7JkxwJdyHTDrWMmqDL6JEoDeaC392Kq3cqR9H0a2aSY9Jo8GRTsEA6jbkeqCWrwyj0tf8fVIYabb
C+S0hRS7CGKTQNpsZwpnoArBu1XYyYmRQDliiY3xfhISg/trMhXSsGNv9UehVcujN+81UEdXADaT
ATjx3zUZSxLtRwEUNfLpFT/1P6uaE2TKfbiBCsdicFjGhcFgW1YpxmMdAkN/9HGswWvQY7akgSGH
OiPNey3O6zG4y0NlQedl5v43ZVAL/8ZDAUWrizEmxeKlWBviG+BauER5i9CP25XWWlKRD/GAb/oi
M6gyYELLLn9DObiCFg/7CUENDVY/dNsVQQaS6gIBCktvgA9fEi3JgBhtDqOvH1+v+mdP73aHk/9Z
IpEIOmZneb4sJZJET/uGVUnkoYNpJ0k5+JF89S1sy2KGzYPq/oKwxOcRuM0tLLLVnh+lIqpKLhK8
B50aCDrZsZ5eEvMp2lDKP3gcOj2NN8MMF0ILHXNcWcIzobd0yI4capuTwZhoNfiTpd1iUShymu6Z
LsyXDq7+gkU+tML7DO2ofZj3VUClhf8ScfoH3/C9QOkz7vDOyyM6lehnSUA9Sl8b5BlmTQKHnXF+
/UI0ihpmwMdM+VX0CeML1Tu0EYVcI4mdeT5kGEhcPsGyQkoZsCBgi3NuX+UjTquQrH/9qD8TRR4D
7NwGsxJ3TIccVZtjIO6K8Z0iV7RQwpqzrYw4fPlAoS+ZG1SZlr3xEnoT2aQUt/tEwRezw9LH4wlw
hlLA+9zDBkZA3P8W+N0r+HWb1ZSbX2in1D94l3G2he3n05WO1Agn1lRv1EXZlaFsqWbKeZnQhtSQ
4dtheDOkgbwuKA8uE6XBiTe9ZBN+AR8aiMOJmUmkdnnAoqk5UNGEEOmetveuuiNgMlLtv5Yc8LOo
IKG+GsD1PtYrnU0UwTLWIJyGoOkF33j9tJwSnju8DjejI2F1Y046LlVahgoIFJqdUzK7SdhGaFCa
uHqKc/84nxOYBZ0RdxqQCqyJqAs7MAcp8Xc13pYcB/xaQgK42QKCz0skF7978ZGcy0aGOnOXpWO9
mQh0X9Jz+LUgsfnjtKgc+s5FtxkUVKd0MadsQldTEiFSBY5pF3A2feE0Dn624ZI3SUnDMZRcsNX9
ijZeT+cWC4vBsZde9TlPU+1f3T2fw7k4ZgwhoISXMusg7vjRmAa8ZHue2J9+azMn8slFJi1fS3cj
EYCKe3OU+mhK5IiFSGR/P5+yZtx05QB3TtvTgjyztXZ5vuXHC+uh0lMN2vLLnXjdFObpUfPvwto1
PMtFmo4VHJ0YjTim5ELoUbb8alsGN2ngFpUQp4Nxw07dQ6DNVtUYhyDXi0icQ9OPZ2tx2cc+La/w
dvUawzgrVKnuXjjCKQU7sO/p2TRm1hmG3YA2xTYW0wHbp/0fqbfpCqnDEK0fvSYOpoaUT1GgwOGW
ysTybP7VqZWDTGACO6zMaEa+ihCuJ1UobG4IRzimC7JOVsdrx1YOxPCBHFrrkkWPPsYltkHeGfhH
CV4xdemofR8Xbu2luwKdVZU0tkRZXrhjNwgABLfOutoqRZf7zymqezfJ7nzuxJZ6n7wuv8Ma5KY3
X5cFzjrQZBx6kieww72jAsxB4QQ5/Y9F7aVWGD/NjOcrnBoesXJrFCec8/ZetK932pIX90keWXnY
GiZbF15lju7aSaZTx7l3QPxfKti7S0zdL6nr7W7T7/VQyCLCjCfK3dRchKi93axy+8jH4Qkogqys
o+Rps4iCNQQ38qMMsHDxJKy34R/0lcBDGm7zKIa/1m6KwMOBUFfjI5NEl/1U+g8fip7yCuKH+S3R
Bo38wl43ytCrTPL5/duDn/qyKe92V3iV0yTaYYRrDMv2PBNDRGBJNdR70GCJ1enRx3IB8BpO4oH5
J/zARBuDxAsebYs2AoJCWzKdZ/KbZzYuBCHF0n2h051ywq8kE1b+uqed94eZ871k4C9SQFgBTG5k
LDQGwGAXhl5+bo5zmIJcXJJeQr2/y/LP73rlrHwhO/azHMzTrHe0ncWt6SU/VLhkOfACK6lU1lyD
lN4gAD/WzmWQNUYYErb1ew12UYmSdhz0YmvIGnPIQUd0XjgCh0GQBhT+KQFav32KssY1LUnVJp1S
1NRAwObfV1g8Y9qyuLHrlL6Xgf+0JUdAvQuQR3LyqEMX1sc47vJzQaDp3qGxYeA4vUwgYFYH8rXT
71gdQYDrpAKwcZKIiIziqVx0djPMD5hEVP+J+96orWUStbk6BeN/Df4dP5A3OjubwyvfqApCb1CY
Pl1yZx3McjEmobu0s6WHQouFVMUDIWXJDk9gCVwrRho8rHQJ6q3YpBaidNVYLLiC9pX/k4VEXZ3u
6vekkEy2uKNZhQWt0BcsjHPVy23g9nSByx/LitlTqK+vehkA1HPrWtF212/6CHyP3bARjcq9YvZ+
t+umMDTvjwKjXkDGRnAfZ30ft5RZQug4Zt0OdxmJ9vr/3khLc4SLuvaYL+/yqEhfOfqNO2HgfdOV
1SMPeCJKYvTNU2lAO++FLisBwH+1NG3bgQ3xu31BS4OHGgjeg5KrozmrOzbMuO4YgJ2pUP2kvOuK
tlEu7M0WKgtGmi5YyyQ/64HX8YwtYEgsZDauE1ohcCuqJlBC/Hc2YsW49GfWLAtpOxjluhThwKdq
IGX0bLFFDoj/7IUsRkKpOWJFo5JTBqYGx8KELNS70eB0HXr8V4Os+IMWQI1P2pP2znI4mpOCk98E
dvJwhp+b7ppv4U+nJmLdTYNROT5MmYfO8wsUnbNAscufpcn3xnEwJEid6ycm35jpXcW14gG+739J
2egXCDYZbxxoiGPA6VrqJO1a/JpOVQB6Kt/cX1YvjDvOmElnJ970RDF2MHDutMNaJuhgSDuvi2zL
+S+628RQwPTk9AbfD2/FR2DD4x31YZADKaxUUIxrbcgSxhpls0Lmg8xQtg51KVSVpFZCYmsHgLKJ
95OfPmYQokBdX3E+k7VtKjrVKppjZcqQn5eaVFTDk2+Oy36udAPuPS0mj5juyS06z/l/0qaz2xsF
8Oe9xp8AL29rMNhLNp2bIxlwA8I1AeBO/ffwFDYDMfxxXCzz81ruX0NlcuA4UO7MXfTerCvXMIzi
2CPks1m/kRpMEHC/CoC7MgF7skoalx9QzZFoAcMVDrprdtncYefQlxbkH94PbW74IlDRA71iNy8A
DLbBSKRkz1y/Rr6HeDK0hyTKON9s8t9ntoXZbSMHyll8r/FoGio0dVksLqdMKeFsiAj1cV0oA6dP
xvPO9pRmHAZehXNDmen63seRookUiMEnTzsKvBr1R0fdritdqjTbelHZfHUr15is4zlA9XUlDTOn
69Kw9zhlVIxJAeFDasq/iT+GxKjsUDS7BLloBwHcN8YdYPYz5oR+S+zNc7TbbUrIVwSDqLDiBm13
2sTID+6YFLxFyE90EYCAPh0dY334EALUQaCHApOf24XJYCwdchBc4A7u1C92em6nH3DJl5sGb7Zz
S0VmZk36931Yr7SfNhXSKi2ss9CioNdbZI+GZymdK9uryxSrcGFLhYy0C37ck0Y6NVH+Va6jAYoo
KsYKxhtdC/I3wUiIJw8ulw0U16E00fzuXcNYKZNsv/S3Gegsf1Wyd+FXb5I9+TQSE56cFhCs9ByS
yj3aSoD0WofdA8rwcq5HaClxyAKhH0ujUALBXwM9NTNDEgxz2xLQY/KfKBLx0cfj0kbuQyRH0E8R
kNrmD3gOumMazF98RiBdRfo/xxz+6z40pm2AWpjhX966anPkmSwbj9PwuiqwHjDlpXiNuNJxdBHe
VuG98xSnXhsurb/jX4W45JyD4Ra+EKcq2LaRwQvtXBjRxeUspN9aVku1bi4jEjLlh1feEFn2GnXW
ovMj40/tXZ1OOzxv60gykYzXuyx/iZFQNWov9x0/t0mGwEKsS4aU8kiDr92LGo1xwHVEP6s90QjV
z4UVa6R+iw/lQTf2uymrW5SFWQrQ0UmgbhoHqofMJdkLbKUj/SMp/O9J8UyGn7Fcez3D7b2YOSdd
ssaXOkey6Uqj3mBR25bvQmWGIHbwx5JGfDIEZB2pnD11aKISfn6O8QPTo45MBar710hGDvXL7c4/
M17cBpOA3qMTLh+MrSsyYSnMpWTzJTBYapLeKq1QP5ocY7GkO4VH6/u8DAezFWU35F18JimAG1FP
DGu2NZpIBdasOfeDk5hswYDeVRIrPe8/YzUDb/vRemsbt7wL+2DswI2z2Is8KcUzfOIV5ozvSoK8
MLy8/SuPw5bPuZ1j4hxuaS7ydPFoJbrls+ar5ebzdLBawUOtr3qj9TORCIdMf1brgj/cGctp2wE3
SzVOenepu3PX9y2AM1V8cqOx8/tiuUQ3NzJ7CzYihcm4L0vJYFDOPxW8rGJPNo3cJQcW4n6ng/sw
DqVueh5HyyEa6Ru4es6NilzHCcdiMwOIiAL3kpUjDyChfQrQu1VW4kbR+h0PKF4MfOQQQMkNl9yl
W3eGoD8Q2bnYpA3R0KYTJbzuB583YBn6iplKlhXwj/0PGjlSa3DyVjNeNjC3stOnQkYrnkA3qWOc
uGP7nVfUUwxT9WEweaIt5Ignd4TfgmZvKTOupj75PAixFXOSJavJ/p+9OgmkBcPvmgTtIDWnfJsU
2ikDZ5F0s1sP5NOzhdNl2Iv/QJkfF7cPeax+WrDuSWRDdM4lyq4m9yP/cMbWh10yIhm4FqJuH99N
oNqT/OavwJEogHvwxZsKCwc+yxCh7UHVD/wWDJcLp+mWaPPmO56A8HyZTYZaFCQHmvhkx5csl5+b
N08FSELjKaHFkfAGVM+SXR5E6b8FsFzI3CJdqk+ebFW/P+u7fWj56twHmEuoy//bVJuelc2gcK8x
cofRaColw0MdAP4KxjBsMWnbNEPTO8WkT9emfqj05ycyA54ZaL92dsFU2Prnk9K54eFNjk5IrQHI
von0nF5EGdzcpklxYyn2ePgSwYSMkuaKZHyxxYCyv3i1svv3xJKLTAWEl3zy9cfbHrqD3bB3XuBU
hwPsZuwOfIqV9n48XQIhlB3afMdiAXefcbqbAK53Q5PfL1e8J+ccRtwcjjqAkRpThLIiMnnzeD1f
qNkRfD+QbSfoYindbqYcRwYoylapH4vt+UENoCk7R5hohXZA8YmOiy7/r04zTSMzOcGSOR0XXG7X
v+5260OJIU9NtkyNAISQ1uuone3lY6eo7ixiBin4uSWgW21bhwN8shn4d9BGk4oOjRcjc8/uFd4G
+7j66q/8NW4qhhZaVBGMzXdHw1FUu4qNA6hGwM30VaYDPf6RRZb3YIbxosZ/Tfoa5OoAOiUW3lFy
iSrV5tbqhWRCIUSC5YEEH3rNkJB1/u0eyas7VFJf8TF68ENurp9RMX3qKASCw+OXk40RK4P16PUj
3CRPWl1VgsJkE/15l31VurajOLwqdxV8C1bnN94NE06SZwWAwnolZsYW3tm8w0Y5Mc5UEeboDrH1
f5Rvpnau1+vlq0sfCw0MdhMJaNaoqCRwT+zU0EoCWeBAzfHWa525WgPXx+pajywgAh5depFh+nqk
Ao5YgaLYxiOY0D9CtIfBSWU4ZGxvvGEF9GchELD9x6DZMCgznNhLYlKP/N2XjTasbySR9CFZkK1m
ILj63szpW+QN6ZbZN6Yet0VYnVzc2TYLUVaMHh0vUnKnPZqBYOlVW6hJrFTkaibe07XLS7TRgDt0
VGrV732TZUo0f/BeKCqaqx1+AtEiGQDD7aUj9lV/QOYZ4kz/kLQuzvCxN1SK38J2jP7e2E3sm+ne
NW5GfBPkzQq0ofBK+DCGtkDpN/a17BHWPgm2szyZxxusZC+248qqm/iAPUFaVyBQOy1aRWyX+H/P
y8EoqWiQ4V5S1KOKBvj8UsoGYpZaYMVdw6Vq96STrqeaCB63IivU09qpfffmiwp6lwLVdGFHrlJc
ZCCaAmiruMDbRD6tiRivg50C9lGnZIZi3ZcrYM3gjpgU8X+iC/cYIafpAAxmTm99ZeAoFx0hyyvr
t5jURu/uul8kmH03FugqrAcr5FIIM1dDsvuv3wQEWxz3hPUlJZDvY2SACl8SxWhbFITUjpqXNjE1
sjNsFdoDdCEuducl6NSsEv/Ebffk8YoUDMglPUXZALR7BcApLcWHLBqoCg4mBUl3m5MTzupcIXx1
tBjqMf9kbNz4uI1ePqqlw6Q6GhDo/B0PtiZJoaFyLfEWKA2c1DUVXMM1n2AgQkz8afXmImSPZlFG
wKooR/FTygXYaKIbnNR5IviGE5DSDC2rhRvHfuJ90A3t/RJXCe8kYR+h9sdZd7Qo3+PJXsDewc06
1KQvYgX8aSYIYUR7acqjHHCueZn/R0X0HgPk1GbATv4BiOx71bFOylnN2bDz0RGNtT9jxZrtYPzp
vn7ebKPijEMI8goiqKTn2JjCzOT25m2kXgZINfY5w3iRDYGeX53syhsKI3TeC7x2SkVJU2aisl6n
2/Tdqv9enVIfLcQER1vCIpIC72MLAsOy2wsnrM+fLidHDVPy0kvTvYF/0qDtOzCEeNw9hTW2UT4n
R+VPVCvugu5KSiItlBjVqgDZKrsT4q0AuzTDInBY9/b+c5szPnN1FLP9Xes+5A9qiLBkaUgkvtqz
yEY3t2CFvsw1+ydKkKvwyZ/mL6Lp/XpcWQurFt3Gelee9sle0whEeJpAkPgMQ1oTOuFn0TTGHit4
N9nXuTrT5XTG/YjGMXyBkWt5O8Y0rbejOOmP+nBuMt7gW+FAP/bzxCQXmN9OCh+t2+L2dg4Wd8ge
6EJROKV3hCG82gwYUAqJ3Bp75HwUoJm2E1ZvwIAkRnT7djb/5fdbn5YhIGnFwjmsUxdVs9TheC5M
dh/ZcsU5MvUcX4OA8KCUrzbLEdO+G+vcI1N2gC1L7QSp6fObd/9iQqOLTMOVsOv6SsPSYMU9K+f9
qElALT4MhNCSTfJ37NbnigIzxpCK2TvPLBVkVSPKjbQv0c74JejG0ViR76rQUBY5TfbQHsK0K/kL
L0j0KtmNXSwFUaWVVwseIqCw91thCLWkp+AG8QDZES96V+4l/GSwMOMg2O3k1N1cuD+gmBnrswcd
9PuCEXlpTLMwwIduXIFTlcIz9WTaTstoA0atluQGZ7iDWdvulhI9OYOUOTA+rLRq4ycsxXxHob43
2K8n4E8W7EL9jTft5a0Ynkz03VRufw33N74rYptqB3MLmPYlCYut2NOuAT38SfJzGAGWoc3xKxK2
mPG60ubFTfY18Lz0peN4eZZSSTUvwAhVhl1KlyzAQMwGTNDHQSMZO+YgCKlp5nuQwiomWXhJh54P
FWtxJp6BNLWZdzKXoUyeiGXrUVWDtuUTA86B5PAGYc7rbvLLfQoM1SUZSWDkxpJGtC8sZ9RxN8sb
WR7him1SSY1KkvTIV3y9vQBgowT7KP7uY8pFcT/s5/QxQL3M0krEmiKXeFQLwPEbLTOyfOxFJPM2
SlKN+zvs6e0umxO2xT7qhKrPluzsnkH/JXvXz1L5xMjShvaADZJI+Qzi76PTPOy6C4TUc6oCzUo3
06jIlwV7JUN5UzTm6xHqqMfJ7HWri+nzUX9cnUZk49shT5Sf26PrZ+K+Z105z7di15WvcEdtme83
G+7JvdJsXyU9j7DTwGX6tUo1s70yBvZYMgojwBz/JH5irM4llimWj7ZwlP618qdR0cTsnWi6tbrd
qyJqlHs0yo5GuC7AgYdrWxbz1BROfJ3gNkF79lyboNyWLrMYhfW4NEKlphckU7JsNbpjeKtOwn9I
xaQkMxOGU0Q1iSE/kEZfqRJRtwxc/c31o7w+1HdoVxQBuxchuSiklP9/F3YZqR7uvzVeaDsogS0s
yEga2pO5nAk7CCN3mMosK4uEj4PQxUbxVCh5WukffDhWe7XPfTy97GA1zjmIzJsmrw6yTX9cCBif
UmtwLKdl4jfLrw+4WFATBUKfzTCFS22BmAf2H+h9S5hm9oRIQQ3jqAinhnJ4gPoS/cbqx2j/W6h7
fN4U5obPfXfsBMqDPswMpNtjLAIc6Zt2dc61PCo9Qvovb+JBIibqm2NBF8CHw4/AqMwNjLyJaYom
G93JbMV390ikBXvVi85K+qiHxOyg4E7ORQU7a/3DjdHLfN0WgS5cd+7070RJkWPIkJS831ET/A7/
Gr5fmTelOmOhvven6bXCfVLviBnCuzGNkQnCgUdZUway0iEjG2ALDTNFDezTP+sckNCEzZ5CbK9f
ee8w81JN+RvlF2QpLpBaJiPfQ9Hsh8bLkUzofkxCnoygNb0TWC9anMCPWQcnOJCswLFAUcp/xGbU
kbDX3TPzuKvBGqhD4HoEgnIy6lpkLUSa8V8BTGZLbi50Wr6BZNC+x0YuEM/mM5dB4/mqjxtVPu6M
dSDQ+2TRLoo7Y+BJ5FHIavEi8zf8o52lc18cxmfHibnyvyo+35ft0SCIfCTh+SAtv68y3WTVBjhA
cF9BNV6qnc4EWUfkpMdBKID4TVvehyLJh1jdcH/1r4rKOxMGBNYueMn/njad/umLG2N/5ernwhsb
ifnA+oQz6yhDumv9QfeYsTjjWub769bHXr1G3jEbC09vrAhLzTdyhGEhKHLQruh1phI/H3aYbnUR
2jcPQcF4tCSyCzH5B8m/Otp9MuuIhv+2FmXRMySbNA3NPE3WEIywnM6jJt8EGpjVChm41sVLAH5Z
42+hE/6DV6lPkXASCXwroNTdDoZBqAZ6TrTlYhJGxfKs+Qwm0hhB0BWNZV8uJ24hM1lhB7Ghkk3W
aa0Uu1r4e2TXFmVP3k2/NhAIdKcWMu+lWc6FgH7ngBs0YI53BTWImSiLfXVjYyCf2YNQTjYqRSM+
75223m8N6LRvAzw7nboAjChJzcFHgNrYdPTGKiRULLkdkEcqdaIvS6EqLkVultzUFnXj38LSSZ2E
3mKiGIRHot4O6Bd35pToRvzKGFBqiakIWtDA//IkXr2UYLNXlMYw4cXiJToKCAFb7PelUMsUyS80
6BK8qBp7df33BJ0PjZTH2sDfjlM6KWRcy2Od1FIqU3xvku8WaI6POfJN34Dfd+hFgIEcJ2RTDhJj
GdHMdveibH9g09afeY2Eo9Hl23P+FViizlNq71dT7g7ONO+oIrdRqwn1/hXkUNesXwH1NqokkgL3
KcE0iYYnUljgzaTRbMI89p43ccFkJmXJWZvoOdwBnh5RCFL7zs4RmLaBVvZIb7xaT3SIX6VemD5e
y115O4BCYhwT1D+iWef14iVOkLsaKXZkPXnfXU8KdhSW9vUCbjREnMHYYQQr3bzwZr4xfDtl/lon
hn7RW0/Dp2LL0NKXcDZPR+Lt+UltYGInUDSkGqoPhZyCgZDe7E+xr1F5jioKTT333gvIkzy8jUUx
wvtMcx1A+sNtUSWQSpDYZkTP/uzSRZWkSkJU5/7iwbArVNUQksMbXBcZu9neAw6bbo9KRbaJJhTK
7llrAcK5LEvvSXx4+XZv6DH+Ln/pxr2ksL/tAVMrw9044NC6GA7ly0OHJFMLG/ib+EcI1lIBjX3X
K45V17VO1y4WXm1yytf9m6Zqub2MIZuYcMQulsuKsp4B6rDjLxDvrjIFYzd0Fz2SLooXXvNxeShZ
V+40BrafwQtDjNcUinrgINad+vzJzRwLdzN3xV7usNAHkTsbmYIHXoBLhqoN2FRWBtY1H1EXOBqg
rF8ee3Z6V7EUTPsc2jP6APYMwbcQZAo1+yxmyq5aoPmvBnSjSmpAu4CvS9vQRDuhLJ7g3RJFpJgj
+3+ErYha0/8HMcX0lecD7XeqTpEiFQaKq1vHgKCtpczkvSs2U2Z+rI1wTMgdbkP/DEErs547Nuff
HfIhV40XHrRTmBm7MRgY5gR19mi2yoB0ogA74Q+iy+DtBfDOmz80EVU1nRZbgPFdsAFIhkuQZOka
iCdt4PQb64WWcGrUShye6wBwu4Lmng+9jbuDco3prLcYASvP53Hfg5jz6Lbg13L1Cx5eVZeo5m0V
KiPk5hEfSr1dRgqeU8wyaAUznzZur0qXO05jwAChZ4it6O7BG8kapbIQhJH7cEU77KBedUx6jM9b
cNlnw5mX+q2kAgtDmTZVRShJPg/9H+UxgoOjBUDmYcwxBMrXcdcx0zwRZBO6KYLUeIVS8+nVDPDx
iQO8V0i20fYqasJD4uoW71javHHxwmUw8dMPCwiF27tAJvIMz3oQ2w5j4zp/b/8Bn3r4neL+LCl+
EIIZjMJCmvwBIdH0yldlUhnRRXnGH1RzyJVM1oh2B1D3MPJnus2uRQBR8elNZuvpqGf24BEEv705
ii5a4LPDCYCJYy75s0amcdJI3CQakoQX4ql+9dgW+fFAzYJpfyfTYf+QUc8i2MU8PfPe7JjNHHwT
VtIbkfqXU+duZJ0zLk5Kta2jVdWV1AK7xZN1Z8nyItpsN9KP5FX44heWXJFPfxmowNTObT2wAPoX
rCxE9eNFo1LYXPgct3Ott6dJcBxhIa+VkYdTVdzSqg4D9NpvzFFXqw68L+LdUHfyWzpfkXpqTzsk
4NVhovNxX4mJerGU5gVHpJeHM+hXSgRV/AyzgkgHWsAbEUqJDhf13lTftzXuSiNcyZz9G+6458rS
HxiikZfeXlAB/q30JUHWCNPuZleMusN10mx3N/bW0z2bqz0VkapqE9rOG1gBIFHLmb5TuFTmjnSj
AO45VRtobuhVroEpjcJntMR8FP36tEj0Q0FDNmf6qIlIqA1cpBhlN7Jg7hkdiIHUM5JOic5GFCXV
Zw91QQSZTMgAZsh5/KcXJ+DaGTXdKp/fdbpCZ7l8MHLp3+zLgGqL65qg0ebXlg0/cGM0UaXBvwva
nCxx3kk88jZSYQUVqdMO9DHoQVHshaARRNgdGWUds1ATshQ73kHPzJwjNjAX+dpCjxNcX4w8l6hy
K4z4xusVuPazs90/Xfq5B4EBXaVkarR9HSkJ4loKdNc93koyts8dreyAmEcvu/CDelw6laMAoE+f
zOVUHAMkSCrQQADr7RkHyqWaQ8Grk+qwUXzlhKcHzp9nZ2pxYopMmJ9GG4DGRMoh3SO23ubKor8y
ZgoDKZvCe6KsATnoAVErlqnku3LdE0YhceXwAqQDSPlr/AqdWxTn6euTEhK870JV4GaWQHEAgWtw
8UWb9fpriWFTWHRTze/dloBXDofvy1xby7s+ic2KesmHNuNnLZJcKYJcCPpcJU+/JKisKxj/zNo6
0RMq9FYZ9aXw5Q/q07rar6masM8CCLCEsFsnUpS9wQzkoUs9yhy4bK0Cr0jB8uXs+luTNbgelqE2
LGQ5MZUG6BTK5Wtt+AKnuzWpeIqCfzFg8OMtb1CRvswhJNaJjgEx+sq4s4oyaSU41ZIs3IOPa7oq
DmuNllkyl9eSnEo8nDewOTpQxJuZlFtrngsEC0RbcDnPxBFzKDYINscKP3BvFAkgJewy8+3Wf9O3
OSc7mcqwoIp9FTKvtExrAXClbn4s8yR4u/UskiFIj5X/iN4/oLV0EWheRRIq+bKzlye01oAJkF+g
ug2JuSXGVmclBjFJWsnHF9fw+zipHDKhuRvnS5lphqA6ihxh+5vVSqWootiQxnrofq1pXa6ZskbJ
2tvJROU/r7ByjZ2mI3GiQUYm+TMfqv8994WDMfsZz5Cg1PfZXU+L5Ed2mry3CAzAuFfiBKBfAx5q
dDSNA/WrP2dPFgUXjJKBKgthVOxoJwisGdsWnKDh7rb3GHE3NxwAncn548chh212URxnN5cDRg1t
e912LyrWIQh6FUBF5moEeWezLybIhUOgXMifEytdhzfx32wnWbhx7xPetqkdbbp3puEvQ13PUsVa
K9UVicxQu8NDCZhLhjQ0L2jHVo0rQU+fev04h0cUMUh8N5ivcRdsL8NLxvJTCfaa/mxj0MD6sx80
FSyNAe7bC87rIDJgw3cfRO45SGLlmGoEXT3XVX4TzDnM0keI+EwPkMFAI1owO/Mi0zAj7sV2TSnr
pMJBx5nUZgbpG3jknLrAwV9eGXx1698DuufED/emy2r0CaLBGVuHEic0NsrRh9eSg6TcDFAz8qmK
WR5QIO24fMbYMqV9bMukrnBBRVbR6ftW2C3IS+ES9Y1hFU0ub2IP7j9ad3bx8LJvp8UNstATwtwQ
PwTWAjh5Tn6Y3GjTCou6s3d5VpcmDXu/4E0kT4YfpthwKNl95WsQeSO26+vlyQedz7fTi9w8Eq7f
yQm8vUikbMPNJ3tUz784ai86nJbtrwz8/mJsb0xlIk69BIAeCxM+NanfEVm/ypdDFN7CiQ1VcElC
nXtUP1tGbka32cblwPjTI2F+vGi28rqwHpusQPZXocHPbLAEg/WI/pQNwgu6rYZ6hbKGlgWli8iR
+W4Ko2hflHKz7kx+gEvEp/Bup/fhvaHwisecrJWdHNRgKf1CawSpza0UKBCNOGYi7pzRs2LO80r0
zfkwCk5PhQJUqPglZNnYujV1VzFmrhalr4i6yTMn5i947rBb1kxX7htk0qyH/amlmnVXnttUPwtD
96+97u/U0DEbLxFgkiOlZyTG6OxXyWG0Mm/y4A0vSfhU7W9oXv+ktFm8eiA/7itNgeS7V6wyKReV
xlBbO4Wmrbam23FJX0mNnKMC1c1VwuGkUiZL4rZRt1qHwJGfPiNYoqlek65wLIio7g9sCOC4Rr0d
QG1q6punQQjmnp5CE1bjyL99UMWNFPMGd4YyqJcWD9BEN6OivRKncWwtY3G1UrrwvzD6eqHLoXw8
EdMOliOcHbzxuYzvjDCoFfnrGXvNOQ+MnUREiUKYzf85xXTXr5yyOpeGEK5FGCAd6l1azmZSLfLp
6fwrf3KST1QrLkG4DqvyeaQb6ADgXWv0YT9TKET01nRc+8OAH30bvraz/R64/xTa5mfTovtX2I+J
vl2j/yhT5rMgvleNmNnzV0CwJu7tuGtnzHFJXdwFKJ5P8oWTk0dVZFtw3RPYGuJkD8+q/Q89Lz0I
ecCHlgIUewIxprQfEHvOq64mKe3MrbJMxVHkZF0UWAeJz31VxhDv7HpcEX9U5Fm13l4uaosAeyG7
B/Yhk8ELTf4Jrp95+SGzBtwr1lQt0R7RybejzKswe79SsO6OI8wxPujkhWZnUmb0OlAkSjqoaucO
h0WZPe8MXMdK9DWzfFeH8EKFsc10C2meDqfhlMuDRNcqweK8CWu3bjyhgaDFxc74rMwFB8WoXj2W
eVX+Km8X1LX+9vybEmQixXFEyCQVqnz+lNtuCEN5RhCDg7GtqpWF8VJXzr1TCVl1pQ3oAAuXfkyH
JZK+dZsvbmJgO7ZqLJ2gr2ol2qFabTneRMiaLzKJD9FOP7BxvupJqrGNRg7RmcZiYMnEQu4lxabX
dxi7IzpsGzoxLcvtwruyl2vs6P+UjKhVBIbBpi4Ao/Oi5vBSqQk0z9CxsAqNmPyx9OtklE1XwrqC
slzstGL2fwrNYkWAEKi3if3yyep5EyTkgqJgqt3dsgmtJv+OgsLG6tQL/7XdUMsusYATeer7n7pr
dPPFQQgY1Gr1IIa34cdUVb9waQLMEGjFcUu3fDgF6V7q4aCYFjBMy+glu3ckJyu3EEkWNtvsqyn7
GMznHWr2EnsMseydhwt76tGHIzBqg2aUYDc6BSTPfjpWzOA7jpY+wC9Hvy37Q8zfJuHvQPI2EzwE
82Sq7XWqG4QqcS3BnjXGSM8XN5K8+QeBrrpRyJCQOVLPsWDvityNoj71hYl9UcwPRo4gd6VDLP2d
fMnC6muGt8dN4xviuvnwyAi2gVJqX4yrRnD+NjoYhHWSeKiw7mq2hcqhcEMWtiPRFl1QCP/Mtf7t
lbutpTTA/4rnmxQexf6j/jZnlLW5ysXvHduUmZorbW3d3VdecHyxKihi2uQNHlnNeLlE3OetqYW2
oNBLRGRnrdVAtxKVK0+Ka2yneVqi0BiF+HJbQ/Ixdafu5FMHNWJKSxFYW/vlScUeKTuVl+gVET8h
Axo1FB2yKbM3BK+Oz3T5Pby9ygAL6o8lVFFVE7neUpy3PvS9uy6dhggwVnaJ+/SDIr2q8BhfclXC
eG2iIyCDmcc0vpbkarDAUbJIJorynzx7/c4LNi/jEM6fk+gj/aUt+gdAeqv4grY8JOlvU1Pt5s57
uaWAbkQXMkJzQLxUjhngpp8wVY9frdaS3dfSJL6xr5BkDtUuqGlpFMbFk9VbPaDs0nEDs/qXkH78
FzEH3yv6luR/MzAhvSnsAHIBrlXxs+WTzbErnMhBRYgfnwv/7fV99sJc7UVIWao5AvSV9B8fx+mB
iFnGnqfKwbEw2DLdMnSiG9DLvwFw6w9nAASCWBr69gOvAvThakI1BVzjjosrecCxHsl75KZ9DtdW
x3Y4u/ZYcrCCW/tkiNYLrULZxyKDzUcG5wRJYAG3yi0tVMsUB1XiwU3mI43NzXew2is2PRFLcRgY
mcl5HOh6gUg5bOyWlnnMujrExQxFMoISyVR0nsmQAqmO7hLYFkATp5BMOu8B50E1EiXLrDunGzOF
ksgnf2R8NXjYaKrOGJ5HhmE+Lj5hrtjbZ3Gkta8YZVUl2HHnLPnhAomosEvPKM+ygDgJE/3GXpoi
9eOs3DBzKzYc6+3V6ViRhZhD3iwpfMhBwkUVfmOyY7KmwkQU5WVJyQ9L8dQ2r4LZcEHP2R7wvq47
oVEudz2tEqP2EPmxlFf/alLOkm3oaUbi7uL0OnLmpCR/GCIKmSI/VPhIUEpE4XiD/rbiWA0fblVi
ca09x2C5yjefqReDAoszOMHJ8Qtju3PXzcjPwK5bHrQd+ityGhPlW+Y1MO5+WYRecUdf9/lMFD0p
2z4VzMdkHLHrGvLtrJKnR4yu/NN+c8xyRLGfTUhXmasZOM2VdZjEAuyM7NosOCKA4TZo8x5OlsPB
/XcNRrPhxQu7qjArnYpXPhCM8r5TbdIwNEHAyXecK3mvW0UNLuNKotKT7BY6ZTY1k33fAzLnqPVr
BJEoCmy9l4V52vWuqji5gZJcl71dFj/woYoVqHtaYu+eP9E3gJzc1eLlKPvL69/F4GwBH0Ri/hRf
gzN8KwoAooKtH6iNK4O8C2N7pGfaYqigAcgfWWAl0Yn6CnFJOicn7swNoBPQ9m/DHpEAlo7v1q0v
M/rHFOuBCibiGVjp8rFkpXw7N461I1YrONFEcLrSfn9qbrsHg9NYvP5E9Z2p4DgYR5YtIhYim2fq
XgFwqh5WfwE9dFN2Gfs4QqyfuQp8hwX/xyq6wij70AnxUWxix0P6Il3y8Sq3aLIXfDNB3lcW6mfP
8aHzhyJweIajX0+TEcFbFYfwOP/UtEcaCp1v1vw6EIQm07kAXNG+rwPcfNvrRBL8gptxbgU4qha1
njKHY2X4j1FdYKWJJWvgBPTJoCobwgs8uAMgP4DrnTaFH7I46DvCt0wVEA6KD1QcHayxAVtOCO3O
ZPQ1xFirItS4WanQcclZigwoZrkZwBRMtUMr3pCZF2fPmj+2CBfyfY7pXkH1zb5luR8BE+qr6uFL
haCTR4b8/bftR0jai70/sf45yLotTunNg3hBlYB219sKlQVqtkmStkGokyMGC7RjhqgQP32x0nle
lC2VuABxefZt0SEEWq3SMf9x8CqUSBKk4KVlHdZCBCC+nwT1MCUcX88WCQRHb598L70V/VBf4blV
CCx2JH0ErXXZka34MHSjGseJQAHWyxPlc5+ENmOeftlEcATtQaW5T1K/0AbQXW4Hwf9yHHqutLzy
A5RWI+GOzr7wNSChcnQQFmE3CWBCf/46cFjxhCyfVrCkmEiEFxpf0rXpIuIP+CNqwosVLQ045p7H
fjanJp/iK5B8fALl4IOHXRW92S2kb4dGXnlevyivwSlxubs70yxSAR643ieGSzeZ/XWimkzBsF87
zH0yIHzuf5WfFTFr27G1t86B+Sf2t66lAvx81+/OqJxeeqZQOzTlDpA7WCCNiDZYtdIOUaVBCdq4
3dINbw4p7ciF+KIdpqP0gAcLfql5ujBnk+qsPn8WbAxHw+/9lbPq5zQLZmxHea1bHi2QvWfQiZ3B
2pldioZj6sebWBmLfts6hy92QY/4WRtTQD1IwBSkg6LSZIhlGuvO/DbPsk6/uRw0gZ1P9hyOdUMb
/jjdsJuljSe3sWVmKeCsCgh+X5zdlXr0YcojjSZwrhMYHTVC+DJlzawT0U+HINVb1PVSZBjeXdUl
PiEUiEKF5BgNs5B9KecbEbC2VdABuPrIn3qknQxjT1IpVPLFb8AxfiilT/8pysggF0rdg2o+o/fD
bcWZLSzyS7jpv192O0JPsEZ/2uqdqe/9gaBmdeOCQ7mXhm8NrL5P0LEMlMHxCGxY6/d4FlE6Kjsp
mdbOm/ZJZvydHZUBsVyP+UATvjnNmK1c9DpMV0ZDR4cgCiZAjabs1pYT6C0i4NpFCA2jdvqsU1Sh
RsHaSPsC+HPniV2C++W94OwZd1f4LH3WJstD5LUlFFekT6R4tGWe2LHQyJZgURlJ0HBfh5pA6FGJ
UaVP6RIQd7aAbyPc69RaBBqc1k0k4mDeJ9FWGvT7GvzjZm9FTI5gLt51vU69RV6eu91R3vJf7EBO
KbfmHYTPf97TVDWcLTkaCCRX7LXfRVLaLOHFUxA9yE1ViYcFbalMo9FopbmQt4/DskyvowD5z/k8
IiA6jabNhiOQuipibB/IXX/8Yi3j0rczdgazzPFstH0RKnEODUKDjCGZ/BjwdFMQBqxabWCj6Oae
IEI5Gl6UW2rt3twbZJwSRHnB3CnqJFipcv3j7Qa2/JkNDyiNZ8m9ToSjfiZWXbYdoTkv2xpz7Eyh
trlUgXG1sqoi1HPnWTrr+EadZv34AvKAAE2aRyKmTDWWDnY5By+LNv7ZsOGMNRJU4nT6afyEkZof
4XATnIKjn3NwUyuk5ZeMccEezetJ87bCnMcANfzTtIuy8XMI5+AR7P7TYcxQSRKcQGA/kMZD7z06
mItXLrsIHjRJAL+rAlbgvxbuhoguo6v9YTlrAH/rTgTB+1kJB9HheG4e0fxKyK5WRZpzmKPD8Jr2
4w+o1VD+FTMywkLJyCD9RqzwveRN/qJxBuK9/I0ONDQeJrAdq3M0XajNvAwYVCZI3zSsJnMLzfcR
KGDmA7Ibd8KFhTqL+M3i92EzwBu2xIJq87X382nQxwvAaQXawmJxKP19JjI4p8ZviEceX5Z4NOXo
HrnjzTGJ0pZZ/GPFG1/ToYhGOBHmU60NqrFYNRlsO/6D6EhwAw3v7rYiUdEkJWgz/PgWoRjfrfIO
Rfxd0BsIgm0K4/pBeZBn2X+gDjLgAXG1P3Jc5/nslib+mo2PJ9TPGomERtn7/vkWNc8nohdQtQNM
8YqNzczElYRVCpQz66RVjCvvlYvS03z2xCAuekDEYlZx6jt1j/c+hh1JsqrVhrkj7tpz07SPsq9S
lCpc8lGL70BmysCnWKkXmqtWy+nv4PkuiMMSovYVGR74aeLOcWeAd/Wzmf+nip+p0HK709Yd1rni
uojiw5OH2HgPePUzg/GhoLonOdFfQfYYkBxmidUN0Q7HLF1pZVKGcBsMIZPQYUfdHtnmY5M2NvBA
x6PaoIRnPTJAlNjvt9pCsNv8ncwdFNXgl/ARnAQ7Odc45UfAv2jCul+gzPey/dk7RGo+YaTVLJct
62v3ohitH9yLSkjj/EgDeRKfK+8u5ktOxecMth3ach39oL/3yVY0GYcAf1I8EPJdPCvoBl84oDjr
ECdBJHftYW0IbKvoHOPmfjjq6NN0FPnVPODk8gSReee6R6Qcz0L9V6CGfc0LSAaO290Qza5w7Uyy
YqYjNwvvlXnrJzGsZB93vWgDKc1MsCUF5oIeKJyOXk7otsj9WyMkJAn2yWfyqUR0SIy0O4/bko7d
tQ+teOZ7lXUxHwMjS7XiMScjdBWB3RNmJTSn/gmv64j2It9QgTsVN0UGv/XfpD2CCEDqpwiBOazQ
WMVQPhvYC6A6reo/v3lrAfBa97nwjOYGvw6KYcv38PuthoPljvJKyxbXq9UogseLK6w0/p1hJ1qN
UmUc7KhC/nkeRaWV+KaiY8OauOqrDgHMPGBpK0V4GfkFlhwYMTmBM1fQKyR7FqF8gLL4LyaY9V6S
/HSrFQGCg3tIyv/0AVI+iVj1gsUEEoL6sweOgYI5XkE5Kwio0rASwboPW/UaJaWUhNs+33nCsDMR
WsU14vCwKTqs3CA8YSnTQaaYmT7jRuUTGivugAmas2eqDt6RpsyPPj6yu6yijx8IAuwKzq2r7H1P
SLbr4h95j860beI169Zg1S7DCNfEg3TiHeuu7zGvoUQE2Ctn+UaMpFE2Vcf8jxckr1YhDhcNSdYr
9plWQDWtqOEVolUyMqPjezqiRZzJfmdKzx8ycvZX4eGmVbT0XdW5nHayXOrXmC9dPw+U7SvRWqIP
pdKMXbsctP3ehQb17n5DFX3Omn8gqvCbQmR6/i+mr9Rgx5Xhl2ktf6JaW3lWpqYOxbdKlNh7s7EG
v7cAIoOP3ynTNK5DEgGd0LYBs6zBoVCu/C/Eb17/TyewzJm7J1+q7ozR3m0qb5Ehx794VaijJAO3
HwxRtKz0yBsB9k53MFWfXB2GNWglnXDwteiUz+yre7p+WWmJLP26T7ZHOHG8/TthRyCgRUt1YRof
PMgWgSKq2Qf+mhp0UT39XbkfEJzx01XNffBYfKIqJsrQPeSFZ55d5kDNM2NIKjkXN9BBmnNR32ZL
BoI4AOrHkXOaz9xD8NXMRrtXvWIaRNeKmElQgblR5D+k65jMBTvQOFBGZ8NQqSNKquBIczX7l8n3
Z9yCUU1xbb/2xawPbjdMtiszHXEFBxc4pMlCtGWKUNxRE3LWAIzSs3PmGjuVR6xqnbQvDF3xvJNT
6/XCKTxir31NzmBpvCqyujmwiSYt0jdvDswdWbHnr4BBqJZbVD4QjMGGN0HsN5hmTi++mind6Aal
BY4sRZJlFi3C2fHYSSDSAz23jMMNvkf/xFkxoyI6uj4cfrW6AwRHN4pnLFOkFmpmCD/yNW9csBOv
no8/QFO8lNJbRiVcJ6EJ2NsS8uzCqP/48euaS2qGZ+Vzf1usNKDBqACNw2TAeOzSjJl3M6CgvS9X
wLTMOMcQQNFWeA5ureU4CFAlWyl369Ak/QdvGyroFb/sqqxsedtIEEfhqkKimgi/8b0iKOLCJYJY
WtVO7LwWHfRhBoKwj3hC5EsWZbDcfQXzl07Qs3o7854GryoBgtyEWJhsxxUMKtmZuVC1xhHE9zKB
qb1sbA4xlM1QJejIAINp5MxyUVod5bmPjeIywCnvjM301S8jwYsHQxR563vBfX32Iq1UEmiCiHh1
86plnhUbCapl4+uMPzOSyOv4WIGvkHh4xSVLLzQ3G3RreIw96hKuCye1AQKiJrLR1pujiFyD2msm
Bt4zSrlEnvxlQv4yZc+7BEK/W7dTZkuwhOIh621B7uNv2FbRwYoZrxuC2A/JgMLKR+slfqp4PqD6
DZ7/P7G9rjO1fYEU9o9t2rdmI4Xg529TopFUfCQstr7WWJOPdz7QVn0Nc6JiQury+eHpNNN3B+Ej
A/+KLRbPivf4Yd3EmgqtcMbphOVsbmBsQ3SDqoFJ7i5RnZePeSoUiQ7zlmCFfQd5KXZs0dYNpzLQ
P9jHlYZhWZnrJ3iaaeDEFzk5GuJXfvRjcbk9qtSFtUK9GRGkzwVD3dgfi4GUiyu8cU7dZyAV2de+
AxcLf8XcOTe6VadZlApwKuhj7C1WC8wVHBfdeiWcyN6/A41rrmQ5sWhzMwmdcSRA9yAwe+AUCn3K
EFfBvtGjuFUB8v/DMYf+tk3B2ystAB7x0vjo4um5BJSYixC2J+uefDnkDAtXhqTiE/egqq6olPeE
NIxgdDQSvkMtk0IizeY7/6xtDuSFE0YRIRt5YCjPsYuvW9+b5yQrr7vHYdWyNlVOxAKwHLfw7adK
6ENvsTfel/JTGLgutUsdFceNv6L1eq/Y0iOkcfmqcacqMFjmc1vESaU4Kb8gqkKyJVtp1m0v9Xxo
7LKbW+pwmzYy4wLPM0YLCO6UNpRZ36fQO27OD/h2bR0N4dHVCcnVSpa20DZXOYdo+nIVANklTlg9
TgBKftAdJEwMx1e40CfGZ0VYXctDH+wjD4Z3dOMiOaHytaYTqFnuWJ+ityGpPc35HYh1PeovHifd
TWGVJP6srobTcknmbf6cCuu6RgxooN38DQAlaT8f6ZSBoi9nKK17HjJT8+WndZaxE+FpSSVt2i62
7F3OKVVrMPNy16F5lUqKQZe1WcZ0+537hubAN38bXkXZct302a65Syx2J8iBnF3QKl1RFzgMeP4+
UcoiF7dkHdi/mHTPkIlht7bEPuH2sZItQZw2vy9sixaM/kZEvmpSlHJArtHmjt8G0A/TVhGcofD1
gDG5yAGAeBlkfj6SiXmy0fbkz4VN7o6TrqY5nCigllcjYV+Hu7JMk+V8EenWgBBkq2bggTFTQk7d
nQUn26Po1jcCfqtBC4YtR9ZivKvOvVJO943yIsdR00f1dBf1zV8q/jcUGh/4WY0Zq9AyeJfs6q2C
mLh/UciJ+y9mOfixGDETIMqUd4Q5sezuMc8USvvI8jqrGSuwEUlafGZQrBi8V79BEsGCA3hdl6kY
smnus/h9vFwYcqPgXL4zdq+PQ9BtDe2nD8Nq6I4iV9j0jGHI88oBTWkep/7d8MEKVYtzGv5aCeqR
UhCAjwt311Cz0EM3W5V2Ad0bIkaZ9sDwkpQwxLvudbj2qtqkelSKoiYgIkqsVnDsKctGa282KWOa
Zxr9Wg90DsWFsxX00f+66xEdE8beo4I0GmtS2Fd78elera0y6UDLACcRrs6UCu4raLlSUhsYkXm1
RBGSMeva6DX8Rg7incah05AlC8AWnjai4weOMj8cresQ0ZssVrZ85pLnbw/+2X/80MO9x3XUwo94
iNLxP2NNy8BHkdnEFqO9xN18B7wpiskn/7E//GHgsNhulFn6oXP1F4PrJ/BgzzdkkPTjC3J/oDa8
4VE8CqU28gZpAPzZkLYiyEAiVFmO+Nrdil/W7u4wfG5IVqI5h/39vbxpIX9IGHz1wgBbJOJpepTa
+5po/nVXtfD0oTYZ5tHya3UO65cl91LWBQIE1rz/PpJO/eSqEIYcU0kXhm/5/VeC/2ASuoDrX52Z
0ebqSz4lerKd/wi6vm+GbglBRWmSrqvtyhwhPiQnjj4DpBcUawTdlvnh/fMG20XGJURz8THHutjL
BrvoeTXvEh/se2tYmMUezutx8drOYiHRXCjpofawxVxkhFEscG9AC6CzQUqCoxu+gGULb8k5qXkv
uPhppa5vQ+Q8iib1dXU9tprx8X2gnLFOHTvV1oCOFhy//afTvF1a4PzDDccrrHGbgLXAa7jdWqCI
S50tdUv+9mzUEsz2zoOJK2taXDkfK1Nv9/jfyZJw+sv0CRJYZe8AcyuGkkgC9xUGmnALWKA8jrNs
gA8hmoTZZM4ZMCDoqjFuqbBByiq5KRk6BUc6OcIaB0Od0fpH7dnT1RYvSqir/iMpjjLuLFTM9bSJ
yL9OTFozQYF9cphSbn6FlOV8djlijrDOOHoPfpI3do0kjn4qswgQVrpa9SAmvlPlsFm9gcouT4Ex
9tAtjqhx9i7D9r4soiBw9XzEnNpw90y2n5MAtTzDlEyS0YNeM4D7KHPmVB4BjDwTRAvSidInHy7n
AMK624kZmrPRx9Q8p0HOuW44LlXaFCNeDSmVz11+OxzgygwJjuph9uApp9AcBgG9eA4w/A7ioVMS
kNXcQzEEKtgpTl14ZAjjEeu9nON9Pyax2vx/8z2uLeDZYlfxC+PNh6S/bPrQfify+oizS5Um7BaM
7Ck6W2rFL8SZDjky8Fh5EA7tQrqbYqU/i5eO8VRVB4au5WI++ZXgGZk4jogu5k14wnAn0EhrsB4+
qqV5ZXy7CZ4LWYDcOmYSppA44KSu4BA5Qidu0tc+cdKFjZ02N+4AfOnTaWAuLhBCLdLeln0FqtdF
y6TL7UyMQxbmxzXqYhjNVicNkrAfV7flqA4ZDZ9bwhgvApbQpX5vX3Xjy3EEPMCrbQGIzk9ky1To
bmASLpaFlN+dlZ5L1JyxA7BpaAXkZDxFQlfPE4s/7+FgFtG1ooMmLdN3tqEUFLxONi+kXUBb8+Gi
ZKQcjs+/YghaHCSwyvDu/WtMzk5ShRy6okTvQcJcN9h0PymNQYveiWTu0JrTpr6HKS40N1EoTT4m
s4tR6KKwy1HIV/paE91XgpUGBHhfcyjfvYf7mgymv0qEvrFcoWR1edjTay5kcFu0Kpm3zrfe++80
BPMyzPXmjUmHTBHiLuK812RSXJLBPUsiUojqAChooOdluikPjj7XQFj0gapkAmqRCObDoftUgUxv
FetQRbhg02KsFyojjpWEC9l2yQSKaicm664U/YVSuQ8up+MlosF2+OzwS2RP6nZ4JlwwsoX4OiyK
ghdElG3mKJfh3W37VxTDkLsdrVI60mwmoeng2aKMSpLFxMi24rf8DGKVk7IU1h+BdrUVBbo4HzJS
A/jdUTNdOjN5Pszv7GG8oMcZbavKz9ObIxcZ7wkHpynO0XY/OhynnCa5iWGk76AF4dVVkA0Q6hRm
xG/cJDUw8sQzEW+fmNQN7hnIyNUQku5KRCEtMb2zsDxPJ46CBqVW74pv1re4MOXgGnpJcWx6840i
uBDmwqecbq0dpWYA9hLnqf5dfWr/Nr1thS9ccFmbOG9sqTwhnX+5FC0JpP5eOSjlyACfUC1hUizF
U/LEPyLs6/Ov/rfromqqH5XWdPhBwWWtHdCyILmkcWhRrWXw83+NkgYVC9vwVO6P6UdSiHA/TWio
UG4AhgjNk72qP7N+GgBMtJ+gewd9/PBtWirpoXpf98YqP86emlol9kkR01YKlwxjfsTrNN84FzQ4
sgpQtZTEmf9TJuURskmhYIcVWTce10xON0vXeHWoasFX2KMU9w2cFm4JK68M8lC+EGgk4YNU0RKs
Fziltjh7v4PcEdzY2SXNx7V69pHeMhQ4HGbVUKANgwmR53lMEEqeXUAw3055Bd9Z7hztqDcJoywl
fX2hJEzR2j0aZDMZMxmFhj/GJ79pNIvig+uxCm0XL2obyG1D9pXlJVImbgQFJ81LS0czhUdTl+Ch
VIN1EirYhpuGsQ3EKnXgbOZTlyJkp51JCpQgRff40pcZWxlcFFmFbmBTEYDaw7GGVTnOk8UwI+rh
vORHRVpU65QXSnrAYaA2416duuWpG4Mw6aYBzEU7Z7o/PHU+c1zV+0Ta6F7TVCsDvQUMiCGlHTlK
v5lHtWbEmggiGK6m5SV39bJmeYepCx77XXamQgX2BcdLqvKRfVNorSxZQkygHZKE4kYm8fKgc3Tp
j3qPrzdJdyS2QE7HihRcsc0dOoT8YrC8ZzHHkekCV0yr233umnS0cCJmZm2Pld43dHqWBW6fP6QJ
P7CrLrHise0YsZ0+PdoVV5FBX4yi2Wzd8/PUcHFKHPH6s1GMhO5rORaCMxQrLnX1dJIMi775laFO
TwNEcK6SNP+7uLi+455oU7CQ/yOEVKFbt0CEdx9EJyVGAB6bkZMTTL2tIbH7QtGnRYgh9FBLtN9U
2+gbRb9c/mxU5tIBmIUDDgQZSSRf1beosfWOd4TR7TMp6IKA8gsv0JbSSwcO4kNRr2HQnVMkakdP
hflWHGBayBRQXNbvCmy0w48rRvI5vjR9W6fzmF+uwCsKHApiS9o5LHxiQEhK4dDyuSSpFQ1TiLQx
sQA/0NshSQ1L0G+VSWtmI1vGWBts6ydO3gPds7jgSARkcLruqRE+LL3aHWSZvX1Xo7Ud5newV2xR
eFtW8sO+jAFYYUBGq3rYo0vpJ4aRSAxUGen4BwFjXXZJbKjZFazgdXGDGCdP++tgxYj9Z94LxXW+
80E3ZMv5CqjfwxA17ln6XPk3MC7e9kS4McZ6UTdReLL0Z410VOcEriG+gQFrSiN4Ii/PUZeXoCUv
PTTBbql5+fvqEIzVlGE1MQUQV8+aHJy/A/9q+WlWageaClpCLGIoaWRctgmmPfOb4QBGnFZN++UQ
F9NVjqpbf/lcCjplUuiKBXdYfQYaBgmX1ntB7iAr34uDsPb30hBCyiFdeNDCmlqTwudQiUhYe1Ji
CxaHTF9RN4BIlgUEOVQgUABeEeI6r47lnCidNbRX8CE2o+/v/hIsMGRaqs2fjO6Zj0xIWxzq8x2B
wk1eg4vvW9Ptu5iLdK3JPyoKo7RgQUCUeCURNiOVLUI1ZlA/UgmXM+acLrc3IBB9kxF/4HQsHbuZ
VWxRxJ2VkZwpR/tcDXw7wQkI5EpL4B5+Tjd8go7PxETLgU/Do+U2iKw+UiRKnxq7vcmxERGrporF
J/d5yFj9RdkBAyuWLZZc/VcFxSmOkYe3yLn3a+FAbvvKVuZlAWs+JUsKhoh/cDOIoXVmNmk2SXgS
15Q3twt5MqyZX5dBf00j8JoNG6JFt9DBu4M5K/R1Egj98hzqO+tXAWEPDfYC/OgpQ5Mq97pCKdee
+UJlpvE3f2HQbDtm+QPU1bGlLhAnwtVk9dI2enuCUw4MWg8GgbQd8L5tqhexXjCqR0+KplSy/J5+
TAo6VxKlcvUaqswIxjOZ0QhUjv2CAagpj5p/VgVWNjjfrLrRKoLzb/Bt41/b4wbLJbB3DPZFi2HE
CYBgSTc5w8qVhMxrhZi/qZ3x74EbWj+4pNg61/PnDQaVqYsysSKS9mQFf8Jnlynt7j2vXP7grQ3s
YneYZ7k3tX2YGJ3S4pMm+BBdrP7FyyIkXMO8kaU18b3Bm2FufPGooIdDHgXtJzClBKkXtKQ3gSSv
nex46XHpH7hLz+9yBXnwPjkQssEKeMjROt5W4zRgjqC/IG2sCa9+Y3W5InCm+/Dus2FWU2c8BUfx
WL/Ic9mDnc/pQKsf8J+34qSnx7kS02hXtBn/gw8YH0Yjsd8RnAliZKNyT1MysxBp3ZljKJMHONfy
TfJjXyNHNK5OKxZKMqq4j0b3ASCDdDpqDSvr+HwEbwvdjzYI/0zMx2J0Flkhad1hNNVIBkHox8us
pXAaNgOsbMTf0he0dHxlvydGPMhm/wbTeWLxjt+ZJdmrllSmu5rvMTpkDKMfMvfpR9Wx+hVB40Ff
/SoN1QIrIe/RmNBL6kSrP+CqctWAmQDzwgnIXLMvVmBakF0UkkNtd4ECJo8F/JjMrR2vLC9pcEbs
+bGt9ul+k7ggCPWfuvoxqa82cMkKM0XmwdVIaU75RwgD96GbxUsdgeLn7aQgorTpskLgJF078jn0
sEvZdCoo/i99Q2DWJ0jWNGBi/AhkToTDCMRudFp3Ws5hAnNVz/Jw/7UutunSIewDeeahwCBKu3Cz
UMdL6AF+pg3sl7ita2dFC5KIzfGxJHCOcaHZy9CyvazcEQQMIh848AOQ02Rnn48YjhvygURJ+/g7
aXW9xoMomYk8flFyEQlEq8ydY3qloeRNx8M5kFMRdSFVSZkrXTCXYS4isJZjcSDss3cchDNoLaw8
25bkGgJKn1ahKRYOwYEFZdE5OGKWQU8tv7g2wWEWPhnvg7lfTjrBAUctsLlrzm7MRhxyuFN/jpfK
sL771S3w5gKKaLKGm58TOWvXH5QX0M1bAAaKQGLbmWlN3viQBtdwrCAlCkYy3nazziRNN8t321pf
EJ8w7X3QA1qges4puxHnZ2b1QNPQkZJRjJBnEDXcOt+mU+j3LD3eI5JPn991PRBzot0pUOjfGh50
skHuw/4eSlCkuofRJE2KCpvaz/JM/PNcY+YYl/Kjch0o4cDDFmHnxkW8hcZdMY67TtYh9MEWDN0n
i2ERcAdeHywpMcnsfDOWvexTz5lJAMY5b3tLRrO/9EzFLnTAlkzNa7m8Y4Y+6Qo4iuLnuWEfR6mt
hiYFMa4XJKo4dXmWjQH+AKEIRx91N2SIlhlzMxFNjDguerVvpqJJu6/i4Sd5SaDFIdOLgWCEg6i5
/WzU3rYyDXD/ZixSlMOVtYFkKv8dO8BGxpDjMCVyRIqA4hk+3iBl1TKn7c0bPt31uhJcKiwBjfDH
WG9z9iAXLkV2ry7SPWYB5SnPxCHTb4cewHGXMlm56n9jZxHaa6IMEXuJ1crHpcAstE9isIvSLVtG
tkXshrRsgY31kOk/HXRwr9ChNV3pL4ZWX1eSctWiorGvNHU0trrQnH67BS+vhDqjqiPG83ulvrW+
86Qgcnw4yEI5RyxUe0baGkVE7CSjOb7j/0nDhdQ8RHdQuVNmps6b+AtVUPwZuvTksjfow4cD+Uh2
5B9V6U9AgVB6ew5C6Sb+QKee5evDS4ferxOS3GuI3cg3hD5II8h8SFeBEkqQc7cMMd6RoTaHv0Nq
+r18mJ+pj7UpFzG2nFyvxk/VguOVI1cxMNJGriT+zOo6XhT2y/G5fq4F9vigr9aSvvVppHiM/4cB
FVxEaDR0OtF/6oEQa8RUXsR/gBXGqY5uRD3JHtvQ8SjAO0hNJM/lUODl08tKmxqUEuVzCMzheOcy
xL3EKZcPm5JWsi8Xe98eepb6/5k+HisQUWL6Au9vY2lGbBGzsM/Mhq2/KXbT1qRkhUtSxym0EPe+
T6R+2nhj4jCe2F8uUMHV5aLtcFSvgfkPGXJPjtHZN9BwiDOge0IPFaYVm+456sBWjf9Y91aPLD91
BLCSEap0IKMESqo0owoRb83gg4niE17xvb4dMgOzYGtCpAk5bn9C38YAZaZaeNR/4OeIMYFnPKhI
x1PEja/d70XWikQd3Q2bytfj5kbwdufBlJFV0kN74GgNsLtSu/RNri0GkefjhhN8J05hg9KA+jnB
iahMZXcbnPOAg2kjDb0yMiNrMHnyb3/dBqQFnxYMUcp60Z+9ckhFqWh8YDdmY04xiMJWTOtTwESu
WBc67T30wYrn/oeRyzBhFzYn/7jlJ8EPe8aEIByoA3KAxJqJSBZCdJzGmzeGEloV4R8rGYxFK58b
QSyOTG5C1AslFKnRAsnWlxpf+m2D35cd54GFqg7c1OddOLvlDbWYsjKo+kC1Fdut0nZCf+MJ/ytP
NbD66Zain8wi8R6QmfdxJ4pKIlANas+t6BOpkVkySzyeju4nc0JFWsAa0OXV8npp8ig7zIxbDwt5
DkMS5FDLP1nld+2jHAcJXbkGw0AVTlgxC66bTPEILRH1gmwFHqBpEXfwIBaJ8MAusXygEYu0qEjv
oOu/oP9dW4BIz/82f8p30C/mhyxeFYs9g2dZyiD+NQQl4rxQS5TWn8z9GxSkECloKiQndPHDz/KY
Wg9KrnRIR/A7gn276NCycrJ6WxWK25or0tAyyfOEhTAsy6KieqTqLHpNF42WIR6p9OHsID90LxWe
IWg5VJR+1a53PrizFbnDHnD9fKPvFvCWE7x/w1EjJq5tc+Tj38DcASCMkK0E/OQgY6n7NV10hGNI
MgMn8PmsSNaPLOrdqCwm4jKlfL8yP1vXlV+MizhF56EMTDwfexrCX+pOxgS9CtB7r6sLsFpA9CAq
8vqWsj985weVWfHHLz2mEDV6q0UQpJebT53159fECDIR7C5uRaLU9sXyvTO6+brpWZ6Qq/r1xvx8
O3Tuq02Sax5Afm3NBttMX3q0QzhMf3GUCmjkDTjH70ao96y/VQQkOqn8nXggj+piBrdGScMYWI2c
7FsAb4D7kzk2LMZt6j42WqxLNXwfAOdUVoORsgEN9gemjS+AM0ZtJhyyeU5VDCtf1+S5Hml/CJVD
04Il2Tw3XFZA4OeaeV1RcGuhAF2xpmBQ9iRXksYY4q1M4uxQcBGBYb1hfRHgHS8xf1gHDnK46wyW
O0tC8rZAI05x+VH0Qejy5ALEt8HtlYTRn1JuQT02//ugWZ9vj/HG8JNy822q642Iu1DhLzPFm1Bc
IHdkL4vHroHJc9fh3iyiOdc1kZN8fvGxAsUouOINM31HIMhwXzqJIETxy5erMxVnhcfglhOQkvpp
5Nia/siZ6zhy7kD5S1UKHDvC8s+TgTvzebYRKu7/wh9q7ctuGB2tYNqASPhPyFg70S1KV7edIsFJ
Rp7BgwUu6rBJrUdFnUdTMSis3qePhohQYAs7IYlqsm+pPMUSQB2uOExx/LMP/ZhZHxQySFww1m9P
hKZ5YfjbE6ueu1lidgjqQjJEfOcuUGgfvt4YU/DYTrYRWY3hiNnTxNFzk57gpTJrfq30NdjmE7Me
nFWvHvsjVKAlZ2JWwrpMZ0aG32V8X8nQ22kMAIo1eWIG8ZX2Wc4QteOsE7BfqP2BcZ8PC0puX/+o
PEtcyU+1IEH/XvIHg5ZI4qmjxqznS+y6gJjZoEiHAoaKULY8LylHt8ZlcQgdnMLUxAgq/pKFhbao
a9sIxZO216SRxGQ45ov9vrVRHpiLytgs7peFZ3EpLHEVusWZYMKV7hZNsWsMHbeT668aNaJkh7JA
3BdyD9Cn17aUvy892dLBWO3+JmR/1rsRhkHh6PMRzMVXZIe6tGyEttWGEVk7iNs2B2eqk92cBTDr
PPVMVlty3YnyFf5Uq5EQ/V3nlmj4Se6geBHrQi/WPi9fFsWg1N7IwqFOnuk8VVdNiVNRPTBcyCaM
FtGpKA5lWcy420joV6Uunfp3qqx6gOsjlu5XNmcGWXbcZ5kQvJoOk6zRAoMwF0o1A9Ui3jzxQGUl
1Oa3h+wQ4XC6UalyeSM8DCM+kWanOTEFRrId/39ZaiTjKun6ylfV0m08t9tPtFMS45y5pXAIJ00K
XvrQOBTPrmPnkqvAdeinfTEHMHPHZUrpHEwxHjPQ37Dm6nvsewtzYW+B+0PSGRDAp3OajWYdLE+Q
Ms+exM3skyvAjbOP2nV/JCi1/p1Y6enLLtLGAKrilT95GDXvPT8d7VkeGh5uiVb1DrrcIkMD7skD
OBHKgeuoQnkaN1Bo+cBuU3U95IWoahTCAKOGcTtuOocU26gv2tPeFKG3f0jPSN9qVLSbxxMaJVfO
0KRxRZcove7gZDmJhrtxGv5UCBLi4uyu64/OZBdY8NRuUffpcdkIrfD1mYKvAwNen0XVvX2zEUuz
gJaCXM9NCxRfkAbBgEmY8uxY135DNOdfm8ErpdUFf9wsObhT3HkJku/Qutg2N+iJdhkIwuGpsnw2
l2cytjvlwhQif5MmiGOu28ECDp6ZvmS6lRPf/aNaeEfYhrCIs4foq95oO+AiMy4xl/jOzNBJAdTO
KoPzpd8GhNfMmEEVVEW9qpqJSIupYCtFHtqY4oX5x7Z70Uqf+e1jcobHzfuyZecglicdQonz0zLC
RyU9dFJ4FiZK/uSHh4vrZmgl7W9jNjjmyYWMrbiTe9lHwxJxLV98AIdzaeEGeggCmTH1Ad5PBTix
iI+rZgWv/lB6s0l2H7+S2ILZuYGeCxv94w6YTLjCuJ1uoQYwUe+fzMnM+q9P2PuUXM5k2NhT2SUh
QUpAti9HJcK4ej9mrheb2QpHYZuMRuxP+PZ1PJb/DQ4Edu8WTyHZ2vB34w1zrGTJG7KH8S4Hur5y
VKZknXoxms8kClWZTIiVMm4s6ZXKvEEiUL1/9orkFuGwIuzyr2aBhiGYL6vcKx5q6NYK9gQTBeGt
cvNYXTaNPhCWlmOvj6aMoHEmjIP4R6oqI7Jn2j+5kVGwLRtOMqlZ+8U4ujCYpI3iKIhUgJVgmwOV
rZLzIvSM6A2x4PVHnoVfv1ByzKfO4fY83LL97aQbanEdEsgD+S/v0FR3M39sZORovlNab8N+DzBl
m8OqHK9HtD3Zl2cQI0fAsa/JEybkyqewiRl6cjPiMg2EVF1z4s3qyKRFcQTjqXZvv6N+3K9YFh6G
J2LO2EoLex2M5air5jgDG6MHaQ8MZdEs5YrGS7yDR1lvwK742Ho+tzG/Q8piob9zHxw2OKleIPBi
YbgWhoFNKbHC8V6/bqyTjYXXEMX/ZooLGN+oJegKEuAKd3cyIxmLFGBHzs1a0dExp5zFnU2WerGi
HBsQH4Hxm3VaVBKg1haA7Gh0fghUrYLdk0CXd+Ha0PJME4YY9XJGal8Xj0Fkjl/K/wlK3eizobsg
27yy7JZ9x4gPyo/TT0t0kYdI6e/C2GbdU8yvQzt9Y55paoFi9IaGtjX+vItj6D1qQFt4yHNK4oHT
4arq8UXsJG2doHWEPRx1DIMeEWK5OHzACNOy3Vk6r3nZn38/y2p2wAfUWPd83o9TV73OvATD9W+e
Ln34wobcgRWCT/XspmXUn0w0R8NzWLzd5889zA7yaiBst8BccWJpiWN840HACx7159uPBwP0q1G2
iyhV60rwXKFVnqy5EoRPY9TkBpL9P7zKsQhskv6Gev9aRJdfrj0Nva2uGJejGXP244sZ3CPDjkph
uZytfPCrj+p/Almwl+pwpo9oRixTroy3Vs8avt45aIwbNCI4RFm9Tpr62DuISdBoD3ZcQwT1+thQ
GNOwJBIgCrpvwBXG6H3N5Z8B9dIRFuhKUPjhYDENNL07Fm8toj8W3DmMTLdwwplLB2U8sKPrPVxN
UGI4MTEUkrlIRsz0CJN5Gb7S3OGIfcvrqIGVeRsnI3I7luZBkintklo00yIWpqdLxA6Slft2jkUo
B+v46Jsf9cZwBrowxwmWxlRrEOVkZ21HZjRCU+hp4OqbHcp1HOmby47k75vRE6wqADV4AFOV1BeD
XkSA48aeFAlTovZM/tjJ91NieT98r34PNaqTbJBPOR8LDKh//bsEx0a2wncb9dGy6NUro9mQMi4U
yuEyubf00PqOTXCtGBBi60HLucrPN5OwkcLPURFUr2OmGPhXX/GCi91GRllMzRzbGSkOAALne8R7
jIu5m+Bl80ICgCzu3ATt2JW3iBj058rvGPy/ksG626IT0Sa16RZCofYswJ/PY5iO+/hsqnz5BICi
JAtveXTO8v+b0PbCl/b32kUChVFRnQlc6b8TVg2z4Gl6koN/hLiPnkEeuLpQKuLT8bW+n/LrN65A
GjJTtmtQj+gQrNAXHiNHPO125VUnkxnBvj42jNRv/Q0gTVyOAVSFn7Obfy3swp9ND+8/zcSIoMT5
Dorbrk8WIFrqxujrfADfAsmal7eAt6qlWT1yFqSzmu4PnR/irTF0kAWX7Yd/GBwvKVv6XPbcKX+C
FGO7eARVVYBYWTTmCeffyk5CzUTrnt44Q6ujniYRKo4YQXluDazSOEvX0KzfQ3HBHW0oM44woc75
me995v7whOfciy5dyPLcD3QphVc0bbY1/BaVuNvXywLcbQcXv2G1sH0ivoM3u0oBIT2rZHEinjXu
Qbm1rdbGvyw0VJrvlHtUiZN+YKrOgvSVE+lwvHFFzzowG8X3Id6faD/LPbSa7y/Ki4xHLs6nRpNZ
jQsaiFjwyo6ROU9PpJ0ExHPFkuX9/bR8Wh6Bd4JtU7rArS6oUpv/tT/75TD240Uih8O01/j6cWyV
LXAFWZbknpY1/sgaq//V8xKCmTjiQNWdxv7DFgKBMavMyaipQTf2n8D0yV/d0N26KeuLvHb5yMe+
7tH1RyV/uY8qSO14t5AU1LBHYu0kR+NtC0TF5vzeiSd0Ka7WstBpBz5b30n7mYX1O0FuhaUJrzJ4
7UVfgw8DibHK7V+BL99xkzJb4zRpfthIfPg+vLkY9GQDGqW5bPLuIi2ap7PsktQ9ht3AoBftoctH
Ymp8EfgOWW2f3XGMHhufqQ0tT+aWNzbGoW84p+3R5RiCzvkSJYypOi5K90kvhwj8kdcAZwt2vLAu
ZWAobVpmwswstpnzs6aIoO1IigXr8+2DA74HQwqunO1+ZyO/4ijuloIolbMyBsFO6+MghlLXCcYM
GrkAL5jox2w1UWcWvNHxSXB8hLzn8FulmPElIq/E3K6vLaZwKL5YlUS4h/Wprd1ztfZp5CrLhx59
59UE4jnv2Ercniq3+SiO4u6WPLychTAOn2WQs1ItRgrTj1ERPc1SsHmNfMZH2uTxb50lP/urdIOa
bOJv6vIdFuMhoABLAoRQqJnEEvHdpBrO92hSYXMFuSX5XePVEIjLQM+tClbt1X78k9yvqvGADkao
VKOmfHquXQoc2BRTwX88IRndIsyL5HTnrbqIOyQbBGkdpMbDNeCiuGS5QOpMlKQSG6liqepIRIEV
I/3Woe8IAShqwyxDWm44a6bM2s/5cMBf4AD63JQ52x1m3arYFeqfpcXgccGg0Fr3FlxtQQiEPQro
mMDvs0vdjtnp/rBzu73r/RLlXoHw0R2Atq7VgOY2tQ1h70cjoSpGnM0sXJLJEW1KSgZ87wMq+xiz
h21gGEIzzJvN8BAS1KVYs5dgD/4bi+HOJnemSh+7wX2BKnnbe8cB3aVbiGc5ULfJvxk2b/vT3DU5
KahrPSPvt47MzPIIS7H3mxwc47zv0xZTyg0FWc6/xiEfr1pcLOER3aa1tCfKcdwR7ZUmTSVglvl8
ZfJRAIT/ArMHcGeXYwr5CXHuW0Aeg6BpPKzQGUb1AnY+lSHk5ImHEZ7Hv+NlO6M5PhWOUv8y1ByY
8ihOLn1J//73CNNeB7U3eLBI7lIwHlCk9rbDrT9ai1KD3tvz1NGyMtiRVit77JuqiEWhg2lBlYDD
A7I+fAvNNkD0IpickOstu4R/CDXr8ikaZ6sRR9UgZBmpgs/Kb69tDCsTOC+2UOQEBQzyrPGU0GNZ
ksU2oTQbyDUUR0mrX8DbrE6I7zQab7Nuyls8A6ZcCt+9d57uQDaFZmwqfp2Mwx3uuGMqHd0xiMcV
q/CXaM7ONSbnAEblP50IKsBwUQsOdhlAHTVFb8Mdt5Mjt4zN+6XZiOOF9AL4/hFXaAAI+KqPdLEp
1wwfEJmynhHipdlNcL6n72O9yFXkxCMUBuK132F8F9BZFnHlZODc3LJu5ztQb5bD/0Td4nwv5Hvz
zj/YfBjDhvHgdWycQ1DNinqCqKj4HHN0xyUz2CF7GvI2Tpbx5col7iq+bc2prpa+AF3O1YWuifHH
m/YOKSXIruvNT/jqTuoBfyNpM8EcRGMLaFR0fnjQKNP3zgDkPkXxv1l1mYdWM7Btb2HiRi+ve6Vh
aXXifm2sHNnMKWFT7+9B+GeeBDOdDvSZ5n2B9S1IAC3xwkgeWEU+hSRdQ7dWxltjMk94R8VniolJ
44Iw1r2LfM4QWJ3m/q+1b0yDUJF8PNLyVbn68aAkryzEQs0OiahO34PeWRFaCKWRy/YEopkwc5u4
JGJ48indhQvIWg91+MVePcQ10FECxlxzSTvDa2i68ICDvN6if4XTPrMMcmalKZHgeMVtY/cJmCDn
J1Z/xTaY81Piore5Sdw0G6awkseZNyDI1CNLHa/7qS9ddvhVJ2WpqmffKMxd0eC6KmQxIzZhHy+H
xKSRZfarEHK323LFLlX0X/77/s2vXtFSzc87NDtD25VZxd5fdaZR331eCCfNkoS44jbnj3exoypv
dxkE5sRwbqgowheeaqEddYBR+PVkYCdebz2mZbhWxjFgDkFkZeA1OyvljVHM16KFHPoCJdcX9cIk
BA60qi024fz8DaclC832BcHBA3LYtBWVd6AHpBPCxsEfirXnJZGEO0eoBBXxo5sGQm3jVTQ6WPto
wEaB8xYRNOIitFhQK9KrTudgYsDQa044YwHDqE6J3Itt7d7B2KJaTHRdNsMfnAE815XHyM+TcjbN
xMdQ2dw2azoutsdlVdYitulyPHkjCU+JcizXJ5F4QY+7T3OPKCUWfhDwi5mZxxLbflSpav9+dewH
hgw+R82S9/78z8RVRqUJ5CKC5oHp2eevrnCHRlb+QgJN7tVBkqaext1bKuB+Hg1N7tr8q35YsYCn
IpoVJLeuEc9BUX3LRpRCfWctz+18J/D2Y4aM0VJrTHlDyTlEYxQp4c0x99Svb+8nPKzmD4zowtLs
dnoY0kgWKq8y4aLMVhRgQtTKNveMTYmfBPYIkQl7XNYPvui9R31DF5N/10gWo9YT8oORD1TVdgXx
hUHUYg2thNDMeOAakHeY5OjX76Smgsylt2TVY6kmhWp7AwDgCD5fY04VihZgD3ihmXWPwXeyJ9c+
gPulCfGJDyQkw009DFftkyabaCXoKm4Djd2dQGjQ8OMi8Xmm6hGgBjWMDzgibv/OxbVxbbg0LXur
XARIeYeuR/WIevFN/hCDsQaFT+4P6q+ZroophXtxYQr4YJNx9rfSMiCRdJjXwrGRyT0gHjNSuh33
1/4msaqWPKonGzKjWfYtWpDtgKjty1mfOk3Z6nC7N+9euDXMIIrGZMfZZgr0yaIzhsuZLy2iaSA8
nCgx53WCx40n+z6AzxWC70O+Iipekzg98wlaEskxnZIEDFnO+4nttlXUeWsemfl2DO37W1hGS3b7
fwOVM4R07U8t8+qDL6ddxYJZh109FxT43ZM52TgI4nnTr27foNviVOyQYQTYjJHa1zmjM/e3wdvH
YaiK1iySX1BR4DneHKfCQyBnH/QXWMlQVAMnP1M2dEW8kIC3hpy1YLyiucY/ZhSrOTuQ53NHL2Hr
HPJsAOWVSaLVInM9NBzgZKS/OYFN2SpXhIcmV5W+qEENNWzlMud/RVbnBg1yheEsgfOyIn+lBxp/
RnIxi2S/MjAMD/VsDOL9bwlILHiHrcfvoIpJxSf+7d7m7l5WpxZtqmsVjpipAi0zv7cVyAkYmDmH
yepuuhSe2WsavA0VJcXWIOawafnp+0E/sjFGJC3znBNib4or8/OUrA63mAgS91P9AAgQxsWYixP3
fmQCj0uSEnbmsFKliod1ZEB5qwgA4xgAq7Ql38bdwrvcRaU7IDwc3qAgNRCtBobxbBUJvrWqnGX5
7HqCi03lUpSXV7y9T2GiYgslGx7jUEjvkRv8EIhY3NC+RT8G7mmd1QCKAhY0549vXYEQMqvt0nd6
onpM2YAe4jA62HaNlA/wXVJuAvVCL5pnnQHgIT45eBMEDNLBq/eFWiVItmXVaJ/8dYxfP2gt51R4
DBwM9D1tH1jw2RZtEIUe5fthoGB88Uurwp5d9iaNkHIq0K6gOb4SmlibSPH+Dm71BoFT/phzIqAz
el8qkwUGRHmb3eScDN1xZKWpDsDqSlNc/LwLSL+JA0BJGiaAQ2gIkNvfTzbMSdSBlHX1xAeqPFdE
v8Q67i2fdKOd8GeXw6+le7rLj30fT9qFw0v90g2nutCMF4SDeO0q3nWW8D4YvqlxNXIOLBz5o6j/
YrW+6xN42j118NDnXV5loO75g+B6k8O52sieHrmpQpnVLnjlCVzcktU2jO+6XOLFTQ7WML3unJgK
y/LmhdMhzZdrO6QQwZJ0o7yakSe4iJHKA0PRfJPumgautypNs8h9z9ZAEol9CSpzJqHeGgAsQmmR
33r/XpFuT0//JEjdqFp9Z6xM9WdUyI6d4O8SGSrgIYBQEGhiU+sqrkOBNqdrBp9mYJzrNqd6nfSp
obTrJvimCAOW8oeeaFkZ7N6iuNxqODGNkQnrLXEZnTU2pfzp1KzTppF8OzX/tOC+KlqgSwnHWIim
7xFowZj924ggerhlD5b/Webfzp/ZmQQ62ENC++cBZN+xMa5syVPU3oHiQF5yTOpeH7ElJgELbjJy
dBYEtblOVf+n8TBO5TWFHz+FGDWuaPln45ubbF0NMCwjhx9KCapoR8UVM5jUENwTQxVFc56VO0vj
bWCh4Ugfu6mxsywvyDzEm2teARZsZeCvzXArnv+Pf8v12a5ANkHNStzRsN1cYSBgtlkYwTWN4j5F
G2/cv7vZw8VLX2DwIMud+a+N0HllUjRW0QE0hycjRzhr2BiX/rBS3X5sL6LhHrIEu0mjANolWfVD
OQxmJPOWCf1Erqn/4/GHOBfDkJI7+z5E+JpLipCaYsboYQPb0hqp9Yxga3SvXlKzRrPAwtlRDrAG
zMFMKKv0F5yDoGxZDKWfsrFFsWS7BdyPQMPzhza85luwob3TuQ/+pPtOWvVQek4FCxsYcDpAv3es
7m1L/9I7oNYbWHXcjqD+EIW/HZK4+585Xj6a8loCfceoFqUnfhjXMlFkbVjCk4MFKIw2U1BaRYZi
TspMu8VNT60oseZvHdKViitIK7JQ14mlnq8+SFIWXwyXhlFAbvK187R6FZHogFQdMNdfEQ89jQQb
ZLlxNeC3QiZhtJ72fAvhUWf6iLLwGQ8SjswFuZvaHtjFhDnmt11ZE+HcC6Do3ZfKG+uYvGc0Vd4q
6KHE0kz9d7SZ5cxbY5YTxDMhvNLGRSUioT6ey4NYHI8+d7rlpjuX9+jH/Qed89pkWhblCu4rXnpT
Ek8H/tOzwTrvLTRQ66awOspNdwUFFzZPOdWO+ak9rIhpBZYK6NLgPm3bymPwv/Tiy5qYC3gyoX45
QHb/0z2xfUac/8rHtT242rO4RLCWqtCiuaXOsg828AWm0fAAtpBW4UDr4pH5WIseOD9UG1INWg9X
feHjuua6QvURaPhJQ3zHzty5xHk86akx3DRpgoQwxQ3PL08zuEpB67BK+zdIsA018HvzUuN3vQ6N
mQxmWGjg8iHpBA1WaziU9EFOY5T/57GtIhps6TE9IMOHpH5KlkVDa+940EJFmOSUvZtNJoIhpHd7
5G9vdKoLBFgelBdbT5CHSWYFZiZFEiWEYZMeRdkGGs2qcQX9ihd8ZxCHS7T7uN7Fc7WuaIDNzXpR
pOMPfeHrOiQZ7xivAjX6VE3hw8ummWN1eZfa6C4ayUvz0OGDdUgt6LZzWKMwIm/9m2a+IW1QYS7B
zO/khe/YuMzvHb7P4/2kZH8gGeCu68gIZAdh2W3EHMsMUOiHE6MINv8bLyjV3eaL9xzlYjZGa96o
HLnSSdeoegrP82t8m93eiRtHd72eyJKC4XSGKt39Pq4o0L/W9g7YZXoZqBLyPG/bIQ2bxWR6OMoZ
EKkBF0cHxj6RCAruI1yU+fEcqG9Lsrwx45lh9/Wvifg/QxPdeeQV93o+L/YfMwr6wG2mwnFjmfLB
gWndcWb7msYCUA+uK9vKYKGuNi4lP9CZ1fa3MBJFnsccFvZ+s6s13U6vpU7/WeYlWbyjmTILgex5
+Fr9a0htUgZk5FgbfP179+buc95X6fb4gijF7Y4UhzmgdGJXYEeQyU9GEj9cvDW1cpPyHVJQaS8y
GtgUwQFCvynUXUWAWT1LDK+CbyFjtWyjyouScGafkH7gT4BTfDIfzRe9OmcSUotd436SjQb0zCAW
PQkhu54k/hwEIHiSXuL/U/cj/RSvG6R3ORWVpQrrCAYgCuyA2+CeEXBK9jOrJGVlmkj16IgxqiWr
10bQ2PHKphMKTN7rw2I7a4LDxfzSTgQMWQnLW3vJHwcoP569yL52D+OzGzlUibMpSbnc9KQ5Xzeq
GhGgLFfJSD2L1T3tUllJfSD8e7ZxIrDG7Q5P/pc1M/MrjqSttV3t5p9iz8VqrTto7m/tJXKKvzjW
21tx8af5PPjX3MDzWg0ZBr3bMVji+RTeVBQ2oKEUNAas+zBZ7OFYiMsosOMDR6kID6cpFgd50ff0
r48n+qOgVVL2+hVrQ8JJnmrq/JpIZchbG4yRP9HUbxq5Uixkw4QZrcps+c1X9FebSYQJ1xmZCMQg
c9visQDcxt5alxfqIWipV0Mi/jJbdDPxGC9biyVO34qXjv0e3fHLAOPTAapf1LValtcS0VbfVIh8
sSfUnAb6e7/GlvlTuXKbPGZETGo/aNKzwvxrQyyZ8tMbVhkNknp9c04KVgt8D/dBe2FZTKBF/X2+
2YgqyQr9QCaxdv8m1mrIXOM85Iv1tIaLSyWWnZeC5N81sCzOnBa2avTDNceFMg5bhOoY3HuqNg7F
3U+3esgn1AZtD95MJzUQg0fLJEhilgttg48kx95wn5gDL/h+LRNoaHlZbuwveMbLYsRSJUTr9vB2
UnOgGRDA74C7D2fZzbtfdItedx4gr8tErnj9IIVAkdTmNxaWpyKyk33YOlgTMU0lKOjRDGDn2TiP
hN3O/VI3rUIlnzqJ29+HdQwZp1Nq74uM08K43YSMdF5TbMNOxJ3BrsCU2AuRpJ62e+NyY9Nq4S8I
GNUeBIoYuNJfDoA0D0VYNSiEAqqCIvEQp7kZNiuG13d6FZdYAdViFG64IjSRujXlv8bG+cAHRRND
yVpdy/7+oqKpPw/ZjuYyUG+Kw3/6Kord/cr23SaMbwD3+Kps1KAlFNw4RY/B53sunH6YqjSScoZk
W8wLSfaqmdwprXE9QDDYXQ6WtbWMmbRNd5+eeBD2XfnX5tedF+cgaHFrVeKLHB8WlyEMUnDRtn9d
B3/a+dkARe4vxSCY6efT21cQuAvtvGeISBV5DbHf3GzDhkW0LpenE1s2aDYBNGOCLbbeP6DDdIez
Ay4VlL0AVqUzBcmj5ysiqGsxWDpOIZGKUIFmrAnN1oepePfPYdWyYOZJmualBv00ResdpAbvPVbe
Iu6rTEfJp0MUpx7vv6J7+pmf5ihmR14G8xQIn0//hoxx19RsMCM29Fz0Hwk5OiQlBhBKRtYhpaNg
oVIoMLdl5XIacno/kffy+MbPG5Xi83wrDimKARhGieAHmcC1TvnLalMsIfmJ0AWhEA7N3Ql3XT8a
M6jDP84tx4JteSpBAofzJHZ9X23XDg9Qu6mxTtJNex/13zFU/F8farxJpfXBhnc+sncMLyXCP04t
3kOfJeTYsuDSCYAkdCkKlO8Yz13TmBE94w37zZKspZfIWGkrkLGN5opXevfuNFsIVc5qbzqFpD+A
zcOQb16xd46bLZLVv5XarxQiRp7w8hOeatatCasjkrig4JETqO6mwWUUJnUXRGOOzrSefQ8CBVqS
sFbJJclN8F7TZjtbKrPxnhSHTc7nSUrGnItBS7zHEadzsK18ad9UiVulw/a5eAQttk2zxg45hJ14
Qs6KRGJE85w2hWVDIFb7MIHxfoER5kWYbZpiWmPcA4OuQKwLYluGs+kbXLrvmF2iKtZKYAHhHUp4
MsGWMPDtizKezO2b7xip96ggo2SFru65sTK/iO1T3n/CVNgafPQIX5IyJ9dmijMKxsrRA3sZ1rJw
kGfBlTXfRaAt5ebQWwjiM1eb6MlKNA2RwUAchfOg1FyzQYJ8F6DO29ctdCsWbxNGUzhruBRn6Ml6
B1z1OvUnUj8H/oYETEyJ1dightDV6ssZTU5XXijW4jnDlHyT7e0rlT+oT/pxxhbm5/mAqvq0xiz9
IX6DSAc/foXcelPJOyTWeGnMICxhfa85vTCstR7hf3qJwch0PjAVRnHQCMMFEKP0MbxY6pRqkbkM
6A4IuzrYQYfh2gYQfVnLMRfNPEdDlK9JQzf1VWQBpNrMNlaWezF/p65PC/SxIEB4ghi9qMb80RWk
L4EZHaOn48MqnWdgoP27VpaEGSernMoRpIOcg4JJo3gsvbthU/kLTjKR0uJNMD0g2KXVfdslgttG
fnDAloiE5MAPvKrYjYV0kIDBQ252KW0OMYrrIaIPUK1gl3jqx9MZG8UXIoyJcbkkTZXzQTYbC3EN
UtciTASzV57+Ej+3u+h9ibssNxQrgVqDXtj25TeLDScaPcWTuKoP4pgMZkFpy2yJCBVhvRKPOUko
7xotndbuV/WxVjSUlSCFKRb+x/bJUmHYwtNaZXxwY0Tf1ShhHq3tntIkwUx2U/7k+/P525l8G2Yz
JmINoPMBB7wfP32kvG2a/PehMOXc6dn3AsdIFIt+lTar3pIOJTro8FQC1maBDrRCAczy1H8E0DcS
0KPwbLDd33+zBUQwGf+y1sr4FIB5WQkSb6OwLKnAei9pQ8XXu5SjmNCKfrDVbCYAqUP1gCqZn2/2
8Gi+VoXSpCX4KHcVdxhq2T3eRmJq14zIfTenz8sqA5SMuxCKE/KDjkfYyINCDz7uA8EGx2/tVbWW
nPSjLFaYQyCzAJfuXb/Wb619Rnl2jXJlc3bpImLc5XHdXaZ/ApBJY179tBx3m52A3G0DG0d4bBQY
yUDeGVXhyoZEPBvcFONN3Sk7gGSB+vyV+SPtup8NJ3wRpBCw4r4he0yjSHmvCwVOyUX3sUvQS9AA
3GVystqq87OujsMif0nyJ9n9zGHszGxYc7DbVdQwhJw7MeDiDE+8oaN63lUtkw34U5BNmiS3uXod
zWfmkRLUb4q0hRZoI0NKzMdIglwAoAMenOFQZKAiWqM6TbX+ZcRlVJwOsHWtd+UwClI5jFPqqhG5
HtUuDGczrLiVGISQS7XW/G+2kh57S4d96ITwG/VSo4TUeXJUK85aoy3dRlvAxCXpebLmy8D4nxHj
yAWDcEDvaUO0GL7Z9XzyQdJXpg7ywEuabF748k1vj9UUORW7SRulTcyn6uWAeT/ro/YrSgrVxuML
ZKeh8ykaJsdy40SuPTKxXzqmSDxEeXVwu+7/7lO0nGd93Oyd/etXmHGJTqVWngqgRyo78Em8jkoj
CvMeoPj6L9gm1YankINnfaeIvNWX/mvp3xTjbVGeLruqb9r5L3l4NlyEHpz9rYzgazxdDnDXl00b
6GW6UFvNK6ELB2mxgIO6d35PTZoz/wTJAsGHyuTWF/juPegvJWzMxtxfW7F7FZoIh7L9KC9SOuew
y2VEyTsrvD90Tc6y71IasEXFIXY9ckvLlQaMue2Bu7aPuOeRJ0+ocx+4/fcOlmIrjdD7D7UZh6lD
UQlSLCozXhy588qdpi0waUt4u2iiC7/fkUfK+nvkSX4W8bf3xV2NDZuyEy/T5tJj7AkMjLp+GuU6
kXb8PpwPqNglWT/3JKdijENoRn2frYb0gGPayMx758olb8VpGmICHqm2N/InDfSCmUcqpW4rqyY8
zIIU1kipsm37doWUxrI2m68dtLLHAUkRgR5vTugzZ2xytKHgqfd7qZHat2CwuDQsiUcBwOgjCZOe
/Ru0B/HMSaGkgXRcKkSl31vuZot7GFMcnP8loFAvqwZg+UsS0RcRRKfbpaLGPWDELYUG5N2MojOF
xzxB/NfhHJvkmBo9jPgkuT/NfDjeIu0ffenvwOvUwyoaZaeTV3yHMNAey1X0J4UJHH3zxNvak79O
KXz0JoFKVs5VHVFu/v7tshaNRgImKSlPe3yaQrH3uLc8go3twI293JP/OECIqyvSdB4uJ74PpyND
/O5s39+asU7ulXLLSi+zyg+O+fm0WtTIHpejqatgyZwW/VDUXNrVd4v31XIAMs1ymj9GwIBk5LwT
P1AxPO6bKLZCL5JLaobsjuWHnntA4nAukiPWPCxfUr93AR1AUEUSJWJy3t8OArmrUc0OAngmADl6
DO0+b5bJxNgLGGy/1LZTzYORgN+lg8U2DVxLOjZugvcXY7E6t33uxq1bxFJKbA6kVZXwRYc21AsM
rV8heliyeLaoOjfuLzwcfYL6zW83hnLzQifZejyjkW3fquO6nyVh5z3h9Nu1mJ6UgW4CpMgl5Xcg
VW9in+8GkbydkpErbo1Ht0hqo6hOdXWjBEVN41MORAxjQrcLNiw8eaOTHGeDUcHp2zI+D2gqzgw8
1Ec2ZQrpPNe4f7e6nNzSb4JinDPLQfpiyruCLT4I8VpYG44BVgo6vX66sJ/bdziUn3ICuXovD+vl
eC/46WMtkioLlAAOwv8Srfg94VoovRRIpvVJMzl7W2ZbcxpHj8WgiOqYSNy1gF9qPmclhY0O3nff
+74KOd7le7s57T6maXgSJS/ZaMU5OwZONDiuAco9bST9TsgnEpGpQfFo6+zmOZqKasTu/4ANU3dT
BNEbrZR1eylEIuFxIZcGccistqales5WC3XXiZqDrg6iGmcenpQojxE8QwRlGh5RnKhyyni02dOW
5ECrlw8aZKkQrdn6YKD3GWdiSfILgjoFYiVfgzPmTzJmob3L6RsA0NTMYIiHtm/+eG+uC+PMax3z
W37JEb+KaSyrWUuJnew81wsa82IERQzQqm25U/l7Mfd7mndDMxe/nisaDEj0nRaNYAfTzeq9NxxZ
SmOJp5uhkC0N70urvruWJrVvagXUMEj1xI4tCDHpYwhovROScANrcNOtbYhybyzTS7nguIG8ETQY
KDUpiZ46Q28uOeQ7S+8Bs5WadttvLpzkAd/lGhx8QuHCgGqmiLQs5KhIoiAzqClPKjfkU/s8iIlQ
ClRvpxXMzKsfhEWZNOY09JJxlOU6CwrQGQXGzTQUndQYEDcKv7SOUdvvFt3bc7bSMC9VQR7UpK00
BlDqnSNgbpnR2y1Wxh95OzxfMpxHKZPKUl8l1ffrsFxVdOsSIz1KtyQ20w96GHZVSNI7sAZqU11N
bc/1kVf7PixN9eeMSRIH8BcztKGJAgYRMdnLY4L62iOqlXAgTLvM91al2dZaTiqT2TiXJP85wIjS
S8togdNUH1Np59rTcZb+T+nkTs4ukpIhmyzwv1+1PRITHXNRY/NAQ6JkllyNnmHh2xfaxJVGzjZs
6qzKUGrfXUdnBIARdObM+CKvsXnrcvNdmltvGqwKOmDH125Iy8121DKSCXDzO4SoBvlOG2IgY+V3
meTiYfD4dKLFpVrqztcDhxU5AN67N1PYWczIKD4dCjT57W3N43NtfYqlxShpoN9DNwo+ZZwQIouE
eCbmuFGIpwAsxejsqKYfgRCxtsplk1OzFvzGb5XwP8aQ15lqNnn6Qlxi9V9FRrh1GICqG5Q7XrwX
7OLkyKhLx1q51XIUHsfIU6hwy5Om9y/OYKnrBLXxTMMbdjxT5759Rc0m4eHnwM55zAGxvjNEudk5
45beWudPR4WVWJYXoF1rh/rHKGL4pSfSKOgS2J2VftMEpaOGPdBkOMoixJi0MuoqLP2EfH4WUbQd
Zdqs2UylVFew0Sf3M01RS9ecPH0PCrO2YcB4WxNBW+nfWOdBAf8CdwWZdg5SKebgFiEGWyA32J5L
1sy52XQ9urRmkKAmXBprrf/Hxmrl3o7dRUSVQrD5NpO+gCvEg4s4OuT8bLhZt7Q4PZ3iEMwefW12
alh9HKN8LLXbkVocPwVRBXI8yH3dKLqxS7nPOH5djuqADYbBL+GYUN3RUkakg0/+he3r19wa6RXr
Ty87RJTrpZF8tgQ5jYHKek7Ue8CcCY6FeLLqZMdbSM1be+dmUPRWycvzLHZQsvGsMX6UQS8UQFm5
UTec007LTTEES/6wWAIR2KX3HwuO6+BYUEwyuVWe//bQVqCoMZI6Oynzfk7WhBS8evgE+qKILPP2
0gZPmaSbznBpemyhp/t91ECYWYna5hogBGEbmpQAVsj3R8hPaYgdM7kVJco6cFesHzR24hYjghjH
TWizQHwQ3TM+kW1AlzkowGG13gmVUAnWjiD0a3a6yzXTThPqb3bJNrLvvnPN0F79c9b3luQ8fCDi
ccMVVZcc46R+lCgG3H5g1ZlsQGMLilqbhkcuiabjo/LfIIy7QsNmLPCKeMbvl6CkcXM0P4p41890
LmGnOyjJZWhTySogKae8IWpXJ/eRxibKBCVrOj+LbUxE1ozSSoTkbTn2TaljGLkRL/MBjt50/68+
9+2nxYNbNZRLQK7IM6bHQ59tNP2LW9fSv2Pni1wZPMC1ajO0kYxT8l2bRb/48HeArbUFyExFxoxP
vACFXGutIleeaXYNX1fNIgDcCDFCG3JpYpxkkjtapB+7H9iijIzKD4yusD/jy54DPqEne6PlgVVK
0FwY9tsqcLhSwCwoZINxEaF9ksrpYPl2wUOu7F88l5FKpZoOOHKOP3GsLq0Wg4bBRd8rR7sFKrPz
kEWEr4q6kDQhtyLAm947w8lvW2Vi69HqgzMYHGSGjL9tyy2gVeEX8mWAfpugbKURxV4nsNRfE00E
h7QJiPIXSyv3MbJ10huyToeZlwsLmYSwo5Znp9UAl4X28xQ4OXyuwhAifz1IwscI4a3T/+p9XhEq
+dtFp5dDbkhNta+AI3pxllT4NaDKyvmMwE/67rgdqjKWc3CSqjxrNLz0tt++rCjHijMkKmwx96Tt
6SC5+w+IcG+kye+K1Kxcz10uXv0sx5ES0bIiWdVoOVt20MEDR9P8uJw48ObOWMvtwWadCow/yKZu
SRhUH9KnkOOlNzV599ZTSYLI9R/nyZ6QKZwyWBJQZGdwY4VM9Cc6DwSYQKvmAAu4yi4pA2960XQW
9m3cgFJTWV9HTDkG/AElYKuvokaH1uB+YZWTsxHKQX4pipelq772o4r0kNt7MN9nwI24qQkRmkUq
DY3iIrZssslzJmhukjOJtdBFD1x7+wFavOD/Bc0jrifxjQM/Z0F8WJS2JCchshobZ7BAimUn5TVV
MM14Me2PQoBhjxISJGHhCSTadngztua7sUahe+tmNbPyK4qC1R7QwmQDPpv/A1O0YKQ7GyuxY7z3
AH0WNIfiOIPXeDFdChyYDJCnSTd7guWL2W2yMatA+BaQsCgj6Yp4RuzUfY7V60vhCoqYRevOxuwi
pE63pHB0QLVKNj22pO1S27LUnsxVHIlZq9dYX7qM6BGj+h1e8XZIo9gvUBHzNZv5zNNS2SWNGXt0
R/s+kpBneMetfuWDdTTXj/qIZmlC+LK+ceFks7yMhR2syZpznwu00JPhfozshTWu5ktmn6yDZELW
LJchcKYa4NAzbpPLKC9JyVbBLdg0ZPC0zEiK54Ngi+BzH8FJ2JOHj7tyN2i8IPFeF1gT94oRhHE8
4CXwG3wSbnkvXop5NOU+PGutXTz2r8v9xySh4vGDFYEXq78GXZJ5p+y8RyTmDyZcQf0s4I/9fogz
pofnEC4SPYy9eDi22tPmL+PH4S4RFSmuixP22C9sRu67SoszvF+X9scn4sgbiSNhuEmBDJw1n6Bu
bmT5w3L1BiX4FqPVW5tXLBZHUMw1jmIK4C6KWUN8r7zPLf9kHmvcZfz7MxJMoY1DiBc8qnwlCTTQ
gi6xwX4N2WOz/v39LPGuhSTn9B9TMBlImsF/YU8JjzykS3CLgEukbo06gWrB3omVd5aBSyJ2offU
1TuQaSk8Fymx3J7N1ZzJ0NLlxrLG25SsKiFF1fgnV+0DnrVl0HdNrKf51igB2SfypPHmYV91N+Qr
tj9fFfi0nSS5w/QDcX450HQbY9shKmE9K1B9kqlccDsHIEnkLdpx+cETEN4eFZpPKX3gcj6L28+/
NCB97oNHHSHe/aOMnesL61KqhGDIgms76tc+xB+AJWq7/7OzSe0YdaKLTO9dn9tjMuhezAwD7wb7
s6J1LGvUdMirWdpToZxH0upmL1nF8ubS/lX0dC/4bBhK+KHO5t4UcuNs1Q1GmSZ7efJUdxQ97YbE
l0uHdbn0oo7eX/d6I1aRbkcqEaJ2LD3j4iHLxUq81RbZ+Lrq2B+mo4Fzp3sryj2n74EoGmduKlnD
qQZOmr/iPsKbhxGRO2I+hR22Pte8GUe535R3hhXIfERW6qYkT5BVTnjGb2tYPlSKhWZYuPZCwOjp
IxnDt6ch4uGfsGnSTAR58f8viYFMtjVFjhlqV10aaH+NkXJdxKswq984/fGP2rifvEYQPosVKSHM
KxMnPRwW4nW/Df3PDx72wIspLWX1cZwn/tG2VQRL1A8aKkiNQFU7flQbiYVwQrsNwNgSIzaogwqS
5GLMA1C78PK6GUawOX2dK7n4xDuE8GKScogMuEBVGhjbBULkGv7XjLzPDErINrcOgOxavGBbDtsj
LuvhME41nSySRCvGCx6DHoWcOlBhDSbgoBPz5J+lhEheuF02ZjU5mcSNyKyyQWOFB4+v6pGjunzr
d/y3VOyuamBoSdT2Kr3rZ5uV4EbxSS4b8j9SinxxMt/L2z3HH8hNXf3CoPqEUKAT0Vv9b3xDUZPC
h0zL0PksX0wIkSDMycq7Jhu6/gFgMIRY6FpKvE6tTDHLAHaBTy5ujNseagskjtobCsEZ8NSb2Hux
+HBQDVmbbBcJaNdGzxKULCYtzp9rlEF57iVoLzxrUSgPZgGQoxhAuprtg1C747ebMggGmxXopKuK
KyvHYWzoQLUEPoLM9dNkdAN5+Wl0H0UWpfFDopf6fVL0nhr5pPggiYJd2qbuA1G6mkYIEyLWFfB1
ltZwCXn1bL3mNHn1WMJYFLMZCqf78o1pyfiujtzYgr84n7QEtHa+cKuQv8XPl3MK7ncD+188FjPm
REWo698tY96Bd0PWQ5ASOXhuTEePnuBoFclIfEoGZlCpG3+52xr5UDtb/6Xig5kFWDU6oftSlYxm
9guc3FY1VrQ/x52dkGQY4ebu4APd4a5zrZCyowVyzOzJXMtEX1I+Cg6QJQpwI1MJ5xMGy42P4Kfp
g8ete8lgO8ctsx2vRotRSEJs5lsg89VecZzLggHCXs4NY2PWDwPsN54yvSJj+UVGrG12XcBqHZIU
XFzSZeUlErB00u1N1fdJNoO9POU8H+nTBEKbjMJ8T7Wd+ERt2FKwpoEaIqnxsUnuM7wTYq9o6RAx
IbssYVxSQFyA8vFARwIph6mtwYzVzyOL4/8M+oLKj+QPyU9uxXO2EKLplM9mKII97myxaiCOyPJu
pRCeWglTrE/2l1+KhSLrZgCkYuNgPmQp8H88ryV5KPp4rMB0UsHfoxdPq07yOz+CwMA6Cg4MmhO0
yikbav0X3TSCfp4oXJnmDIxRS3BXzAeYkapGG7qAMP23bE3ZCRjSYGds/mprhUUTiwPKt8QEnyjx
F1PHs2BPPl3ndhdAyxIgzlFjpugXJ/c2fnP0E6a13EWnLdslOJsDKm9+FNdqSNC3pPdJxRPEiVl+
IfaGYVHAjd9PXdlpnlXsbxHgj0hKZIvh3OcdegFyV26mHnAccGNBbpKo5wGmslTlKXXskf2KnvJ/
m26FJUj8/7EBVFXrnJ5EmhMPS+hIFFso85QglceY9BmgobtLXiWDdyXCug35jNbQxiQop/af/8F0
JAtCpJybwKoX/e3x13lLEz5CMy5UG3mrTRWPEbM7febjRL+8uw47KOrq1RTDxabI+omhTBE0XvaA
ayKtzDEXi8WfqE2Gbz7YiWzhW64vGxkfbDS5Y4VvfjBOK5ShvPuY6f+uVUWpXryFYxxQavTqI5dD
TUwCQ/bJ8LOvMbf2roQgfiOXtHqd2zSUvyiXbGvdPrZgxj4BFcD67TqEemFyijtssdtdVD5Bcxwl
BYduxKqaHUA0VO2ZWHqPITrffb4Drcdw31m/Ce1CTRP2foZtqe0WfQ0RP09y1MC9xTG2dr+ejuNL
muYIDMh7xMy9d6HPb1BYPKThLgOoSKqgl1TFHyUWT9eLmMxCrhQ2iZEEq4lYqGEhVjCoq12hx8DL
MvgKRyJu9PI5F12N13jC+8WjtKfk0+2wuw1jwfxN7stIoKIs9kgGPGylNhpUSv3BpXyIsWKnJg8X
EbZedS6Q9PpWGua19c2ORqNgbh1jxDOekyUfdByg+6oAOfnLwfdpuS6WwDgaqygxyLNdJXHorxPW
f8v0ZF0nv7FU7qnQJqSV1R29vz/k2E5D+u9jrtqYYTg3HquzA49LEFRHmmwHuQAqYup1LEg7eh2B
dQrdExRvyQ/53BtKTz+fQa2sRN6AOzQNcOWaiygCCgqZkn5VfKPr2P1i5m5KTfULRmouB7hsXX4m
EQHZDuhrPHnKC51EYkk5BkUR/IJnDkSXY8lFUioSAeXX/CLzUJ6XHuyquG2+zhU0lFdOtanf3gDt
XSRaoUsJ6McI40oEw7mYxn+hkcl4kzwGPIpNCz2m3NF6NcuUyZk40KnI5g/FLXNC98dVZWVWbrCG
5g3Czz2u7wJPDb0g4DCXAiLQ0DllEGJ2eQbKk4ENqc20EXJEmjilKzEYXl+qKPF+4ADZafZ075gc
1WmKc8tqPgwKSBfRv2MHB5WVyPANPZNhlaSAukjyOHqA5HJHSHxgBkK/e67ejirnUMpGrV9pQHln
PH+qa4M2xhEaHN0AaU8h6hEWWZnquVl72uO1wYTI7e+JVvHWa78hejNBpXF/t3gVaEiRobqjFRRK
XI0mBjtNRx+lByib8UhGdjy+G0k9ATJSEVUVCtGdBAFMeVUdk7LJdAqLXuRkIqUfIO0Bfj5VlBM+
caVGzesSGft6A2pALIYi6HqyZ4tPgW7+g6ZqVNeHJDa7PdPfSh89CX6uOzklxMl55WODbH6hg9ct
8rUiUQigp6gh1QDECQtw5Wy8+IWDEjMOKoIhdfsrf68QuRiskH+IZ/2ZKDAJr02l9Xz7rqSY2I8g
GP2gFBQvikBJpxb6PXXIGJRSQJ3MydlmHBzNl5goLQXNRUUN7B1EY2LBZzhTxKlzWdwFhS9rji1o
6dGesHStAh2iZQGXdjKoIe++eodbicJIEqmxqoyiGF6r3AYQSMZ8c5uutIOpFWvHny/F2EGSfSvK
mAN2FxEdxpvH6XBxecz2+CT+AtGDnUYeFz3QdsH7EjjjkK1GmMyx45qOm1It/pcvupkdGoxojrdO
dzSCqS/Dei+ftYB3nO9eh2ebwKlQ4PCkPro4oDqPuRm1lg33IzmR4A4njoDGKeQ/Yiq7doGBnGPK
7XZDlWv/rCA4A9YFTl/SVNaKYcjW9VX3bP3svI1OJlxOc9rcCDXPgBzQtwVV3/cKY60RDb4T/yWD
/Qrv7a6npME55IfIDnqwyHoAxHI7sbECECoHg46w8FLWajlWbasXE2duTJYNKhL38ToTwvzwwofQ
D3tqWsXxskIM8auvGHO1nQliXZtt3Hjg3zrEIrQIRiKsA0PqbgUAUbiA/FnNQV4Elbm7L9NVfC8C
MDr2vlO69KJHvEJPc/NTjtPpKDCGsGJr+vEz/fOE/wz0a+0InNMcP9V5+lUqCrY8xpHJ174aT7G0
4hNk3ogwnKprjMJpXtDfPJAs2vbnIQ4JfkDEJvjdpUfbv6tE+G6NljgVdWNSFZ9MXwSWpqlorjew
uqQIqrXHECxQoOCLg+rOnIbhr5C5KBYuTR3FmixUqGeAoxQGMxtzonDtY2+0Rz8m4lgueneNn67m
U+zfLEYi1UP+1xEg0kwDVzI9nhTPVLkNLXrQtzO7EQVT1X5lQqvGDK2A5YsGMrBEs2SqPy9uYjon
fPR5SRoqHMwLmLGv+yoagVBoYuozUvxrpGOn3N73kpb+rAPaJabRkbrt2ocOsiO5t9PLcB+Sn/fm
KbuY49PbnKiH8wcDOoD4CNjfKWI2jieajIzuW+7pkUNM2ldOVsXtWxmiTu4ip2H2QJ7hnPKgWW5I
pUK6o35yWOV9iaE6VKluCHJJ6iLx1JCOoZfCb+N7YPt9NSKNTLwwLWI4y6akEW2nCelILbph4Nhv
NrS8aTtgeUOEADv6Ey3QJqqpp3ILeaTsb8T9Khbqd6CAMeg6FuWN5zixg1OHf02fvlZk85A26EPD
qbq5N8fkjcH0064zq+FwjmsV6YUkSikDOffP6RSMDpIxMDEXMbHOQlSlcbs6FQYDL+9sxmhkwzuv
pULvsn/wvClDdzYpJD5ggToZOoaJBovFYCOHdCxBLzNunHkoHcMwOcnu7sXLXAbKP+x9VJ5xk8LC
sG2YtdvdfCutedkCgCmL7DFlrTloyxMnPZ8ui0sRogOQvy5miDoiDNNblOG3XI1D6w/Y3rfbiVSr
il5h4Y4SYvKgQqKMi4I1OjIZ9zValbwq0ZhAg2EhdcJYghXhASDLfxofn3FhSExI7D5XUHTlWDzZ
Rykvsilw3TzO8OYjT5JgHpY1VPYk0HwLV8vH7/To4L/bnOaoXC2/zDalbZBiHSLqdJJGL6FI/2ar
otUho/OT1Fl9toKwNy9Wl6/HfaFWbZ7XK9iCT/94dFF5YykjlWdXIOZ9D2+Op0B/Umf0jsI1WvZL
o76fymdFLOceBwPodxth5xvNL1lc3395SHHm6h7CKhT9NwFJPDfflDDcHFnObMlQ3gP+RBW5xIMo
2A899qMuDUAuIbxs0N0r7NwuaHCputBuR7EHw1O1XcNnJ1B1MPFw9jnNPDWki6B3IRZk4xea5NHR
QCOPkdjqmUs6NZMLYbDDE9Tu4YQs7eqVyuxxGUPclD6TjtT/bamC/nEDde+w/iFmndcfCkBTbikV
ZTfRKaesdXjnoTZnCo7P+rbtQpej7njEukIzkDMtqrqVmY9Vgut7Os9lUY63VlN5wdaeaNZdEKdD
PBj1IVZVzmdzGoc6y3AK81ajanM32cARdwoeYTpCgnExQLH4ced0hvIIEuax7MsONm2CgZfLHCrl
iaIhS1fU1L6wy4dR592nQuo/R8AG17F+nBmU3K+boc6rwOhDbTFvmLQdZy2p0ZeMQChwvB912iP2
cGirRkMe+jsSa1c4/UmnjALTvgR7MS8fvKBm6R0ajGPxNut7+sNgVXJBWn9VGWU9oyfTvZMNZTgk
ZulDtez0tr4imnweItbyTTmNkw3ayVwJXxkJEtVGea2dIgDAbvJIckAGWOcIXm5ql5Ed3h62POd3
hldVIHElvA/zAgozChveeD9eK3ajBt9S8tqsdFarueUAwuPABZYpGQDeS+GwwBmkCttjrB2WnF+D
xXb8ZmI3aSouGq4BPKyXWwDP1Qxwn8B3TFA5CsAjxyKLqXdd2Klo//ykGCPl0tqCU2hRdd3pqfsp
YXPEf4/QEn6PW2H9EgfHJt41Y34E/FRHB7hWYGjFE79nIRV/BEIDqAHppMsyrgyY4lQefzqBZHQP
tkFy3zsH/xvQMdpoIa3gX3DkxS/RvaCnMZ7GjT9IGuzdl9PzjLsrMn3vzjfNnMylgCgfgLXSPe0Q
LK/4cZdmTbw2hRaug/F1tPP8+prBNX3bUHQ5d7ehOAoeW4dMVny2s5vo9RDBgP/LuwVoPUATdJ7I
rhclGJc95Cqb4EFlh5JMUHBC9hWVjUPjEla9f4i5IRlx10OlB7v4B30zkgY3jIrf1ME3h22Mn481
2Dh6CFHbzc60OuuaWUt/WDplC4NFA3bBQwBy2CCG5e57yj0C4oD5QQN2S1wQU/X3o8u8HTc53kbH
wknD5NAwVIqix/3RoCM8ne5njHZOVbzOQ5UhVWo+tO5Rk/xW139NaGIOOlV4cAMk2JfvvVDTDac4
Gggilg/EDSa1aSSNkThJgr6acPOcveSihJLg65UDgf81wejbgScX3UZXf+V5JrGvDfg3g8WmybcM
gX9+i1/WVJdirKkfD0wMLl7omVOQwtFv0GyqFrizu6INszdgM3hJinGThMDR54oYvFtdTnowJi5E
okUnW5V7DhMC+q1D0zVrZeXDU7SpxgfGhx9eAWC6KdPwxUyIc36hn2cepA81RoWYD8lkIUn0wU/m
UeSkVe0zqgESlaF63iOqd7LKw4PlF3pluy10gL4360kwEU2pi8dLjwkne5kY9pZa3ZyI/00VP4ui
OUcE+BdVfIRCs0Z86BZlTZvvpBfztCxpjc23tzckF7gLbQ8RliUEwyB9WDSyeubd3DEJc6SWZNf/
AulA19wb7vV0TyHYZH1X2v2I0UWebOOWFh5PwRT5uI08SsjdYhTlnk/FmNwADAAHqGbv/D4R+QgA
rtxVs6iNvqcVFGkG//VvzRFpalsvUFfZzqWoN1LvtY7Bi2Uch4OqbP97/igje7wo7UYIRuifGH7h
qs3iv9Eu5o4TTqYAEx7krBKAP6FVDzbGInRwiCnuOXs4stWlaPxTTPYkzm7vZVvGfYEgC7IfIZNT
roevMMg+Nhoc1h9u7Cqt3zW4lzsXBTniL9EqnjOIA5MOfpsImjGgAOJUzcw9giaQcs042dh5bFgM
JXarlx/oeMqQfovhdQcdx8LQ2zUbzUjsXwkCTVngKrQJJeSzep1QLJTWsF92+WThv7pdc9Vyjb1e
RnwQJJsimMZwzRcQJFxdrospSoUPl5xuM2d57oe2bhJ3ql8QFTBosOw096yh6vDe85gzOhhAR6w0
8RRKwAEKB479ATqrcpRxf5m9Drd751CgQIAv9/jCxmhrwMjFhZPT2X7PAhB7fE95T6Pos1l8xCol
qSoj2qO2PFChTK1sOsZ8MAmsPeT0iPcY50Bw1waAUeE70PcxOKWD4/cA3/nwFwuxxG47F1wOdY4S
UPrTD1+DtNIGAETn0ClBDfy70I91+7dgMicYvbuUCNEfndCFrLZnx/dxzQHEyIeXccjdoGz/xIIl
4CPxEpVlicJu0yixDNTF6SrnbbzIsVWruE7sv51/36AIrnKUr3O0suqN28E7vbteThBd0X7ML1vt
XcfRj9Rm1aVQavJUuFvP/idJLIlLowrIfhs6x9AgCvcKwVq2g19UPvBP9lRcSJXNLjbiTy+KusoL
vP6vKovzKLZpeemUF5y87geACrtPkg3Ij5HbpwGmvBMI9PKJao/igRZImb5bM3epV457R3tmy840
URzQGR3254FGBZqQOuJMIJ8fNWw/mPo9eIaKKepJcqNyaCpg+MX6ZLjTNwGncaByKD8TurB2EzF0
THcQhpJADLCerzEu/I5lS0et2PoZdHU3P5K37WwXhpcWxbbirFGJ6qtbzv/Xw/DamXb2H8JnOFFg
oFHkvmRdiYyoPvo+GcX2ZmTQ4wO6NqFkclxErwyfZJAodT9cFvZzIQM/TMhwgZfmJgBNehAhq//U
km17+uQ3DWWrKOrWNxoQHZupYq3CoWJeY5hL5mr1H10XVbC7RKdv1RYsmg4zECE67gZotExqmikE
2uZ2xFsFUkt40uDDhpvVCufM+AYfkVkF6ibLVU5pVD54tn14yEVCE1AlKlkrPV3VeosicIRSO9FK
BA7WT1einiu5oEyx6koh4KcR9p3Qt2hBayiY17YSXTC3B9/4RIScrtx1SeigYBfxc9EOWv4CI/cy
iIxleJhzIMwZLY5t3qh4EPXxbJTrOpEs+CrcBRLIhX/Hrjg8VHz7d0FBp9Q/TLAFlk6ZWJevVeEg
6Wp2QZxQ2sCm+nRSqzRSW2o1E7Gqt0sKJNSLM+PRR1Ufz2k0k2MobQnfnqpHK9wM+3JJl9+IKP7q
mkk6pr6BjYwOniH5NomvIrsn7OF2CX+uqyhxSpUNsxvy1/Sb13xdIia04DLVo2Wj8aiUU7COG7an
PdzHIhR4SrA3r17di6K0XtR+3KGcIGG6rezCDrILiZ3S60hm31QW9b3K+xzllWu7kRnL9HxbcKak
wvmnxMYyQlwgf236foc8VkrAPqjjIhCDQrk80n1OVNVAw7/FAOsxdLGFG2oeVcJd9jmlWwMRgs5U
e0V9xQSVu9LNJqEQHfYBz2v2IUSErOv5E3/ysCXvshSkds5MlLHPzDn/7NR/4rIcTL3oRfvBejcN
N3ETgUMMr3hCzqA/d9brQcWIfwF8xr+VQD5zsrbGkQgyLgLUHbwU9+v3jLVk4Li3vzTrPNv/deMl
fjTEuJ+kPUb9dlzANxWWZ51B9C+gdHpSQ3p+H0DtMDTB1Jle5DZI5HimjF8wZOeNfSTcHpOnUO6q
tFGoIgEA7h0DhH39c5o3ktxIpeHHC5937ZM5yK9NE2gDi6SRP3EWmOGJmoqht+39YvMiQiffknxb
6v2kf46qeUEBnxbqxEjU9L49COAxUigxuyZIXGOotOvQdGV3JPV3GpiIAZIcyPQkl9Fp/bnB0ih6
StCvq/wQkAK5oZdrlQ4pV1ocv8jSU3XpRbI4QNu0Be1rmjF+DGC+YNCwOH5pD3rxIwIhRkEt1ZoK
Uj5tGOic3AgGZObn933rMbwJYS6C9tLz4F+zg9q4v5en9C1ZSxifTDev/rMYd3fI920P+JOzbN1q
loV88eTycBGKg/wlojFyMMu+BfoBqloKpADXREoqLzsqqLdLXzKduGUdm6NqwRqaxSzGrXYSpyw6
QIqEeGU/+jCxiXQnO5sKNlu6/H8/e9Mw6XInpSVs+Wm9Nu9FluMsMqOcclNMKUeepeNViUX1obqK
vTRIubiyY7+KxN/jRlYgd3wKMiZvrVwWkXhNQeV+zaY+3XMjaw1svSS0ztt8Wqv7TwA9FXj5M6BG
NnLKAauKiYzk4yzbGTotlSp2pdqXE1pF9w8aRrBqSnOX6C9aLC1UAJO4TIn5I7pJnP38TuV+aWk5
VK89A3Uw1JT2KwD7VlJqikyq+nDMGFeFs8VF4OmzHFvkwuViZ1ryuIZxHMF/lL6Z/c0r8WsgHZHd
1jjT+Wyazw7W3x1DN1z7Q3p2IhKimM0z5oxyZJZcn6v3/gGIZ5/VrbcgYQRm2/wUFvkm6TCsnHGU
L84vSFTzOZtyJFdZfqFp0AaOwL3Jg1E542EJ8McyRPiJEcpD2eBzA/qN3vQR07xubTKAZbjwpn1/
6xwaaH6WRwnDOELkJ7UH662VlR1uJ3Pq4vh+qG0Au9jkXFFi6QsYkNe6/lgNYr4zV92IDa8bSyUE
vBiq04LRBqME5mLrvwUqrt0Q6C6eW7yMyZUNxBwemUkFURnqWmP+dtw9BSpxE8lgBIk/aAiHfOam
tdXX5ksVABOPe4xXMY5yNsC2uz6zxYdbh0A0lmhkvctTgswdwovulWjPz0yBT+pJvHERBfmnOlVB
ABitKNJlFgAcKkIE8RN2XfiSfF81gHgASsYpmeEJFZvnjAabA2+jVcYtmw9p5tqE7DZ+gI3z6dSS
6kevyCd0SNR0Rk61zozfYMrg5GGE4dwbE+ti9IJPP0YE4v2Hx4inT6x5KZ+W2aT5XZfiTUzMhUst
Vh9wdOyY+mAmjjS9ONv0umYuyfu2VDMW72gQUae1TdrTArnwbhVrLt2JHOm53J/4LduHbMsxbVdz
V2joHKjIhUfw8yQu/iAWZsK3sxAxhiR1+Cn2Uw5Y2oZFsUNhOlISvxJGgLQSmmJMKo+R1pN1bfqc
zEKlzUOc5Lh/n7quoQqkF3XN60yniHzEWwCuVKkVcHRTnKjW9QLsRRqlD7vAnXmUmawKj1dFt4gO
CgXztHDVOoLlhU+PWMuUX3MIPI2pZbg3tkFvRwDj4n7wyBnRlb1PRw+HjfgEh5AA+8SWMPZlal5p
7GqR1D06ZvMoIfJUzXUydF++qGgKYRZ3s/RoaTBk85QL1Z1uhxOy94UmVohCrdYXYcszj1UOvYrQ
2P7BdZwCHU+//Xv3WtGBbneLxxvETKZPl9kCxQjpNkAtwCr+KMU6wiKr+ZDu0U+PGb//CkK5LO0X
uqTqr2aLh7AL5Xnm7qQw0sSGyZ2jPjGrUGaY1JNhiyBRxiU38WoTWjhmkpEHaLuQ0yE5LhH3tdWV
HF1IiA8QuaH4oQU0RB8RQqZO4MZh9rbi/mL8OVeeQv/j6UUMkqDSNzeovS6NmcaChF7BCd82zn3n
z2TXQ3zlr3K28QrCVHw5ahswCwTAZB+lLgJ9wUcosZcouOsmuX85UsN4z9Um4SlpdTUOnaKrNeuk
tABo0/0XfeJWJrd5Tyg6mV19RQqkKwygy+JbdveY1Jpy+/bc//3DmP4CHIOC3L1/mLPnHSvH8Y71
BlebCddX0aeTzxKDbTIuCjL67OOs5gLNFCyQM3KC6WAMBRl3RJGq52F5v0OgXSpMHUQr/N2Mfnvz
7KLjf+KBfzvatuIA5eQNzGWZ0qYBBtvNL7QWiFWwl0twhsCjjBz48s31akSkHypVYc5nQllvrqnh
4N/5UJHNEnViknU/Rm6aKpyIdYpGT0bGeXgb1YhqkuNYBfRB/41nbHYJeyVEDvVuZAAJMqQZAurA
TAO96X1cXRQLkQA3SbyTM5sSB6KtEkCKVMGgfmv/qIGgiUjLt9O2+9Nqo0yk6lXbeyOSSO8hnQRM
IGYF+1Tp+nn3z/IQdQVsr2D+PDQBp0KmfzollsvMssg6Zu/L9ndvEhypMPhnGM7tyAu9VZNzfaku
At9Siz0zApeAXParpI9baTTGZ+SrZ4u5QNJWi7N61GInES2Fvy88v0hOeL2paXRzAe9xRmUh4SLa
k6JljvHQJr+fY6UgBBX84SZilm8w9ngz8+wsgltba+R3onPf9/1IvMc4YHBJ9FjzkWYvqmTe7guv
SwCtUpHPnOEA0d2rU+2JTY9X5v71UzSstQOFLTrc7XW9bZce3DiWlMb0JAj9zlne5Xje68EgOhGw
YaatDbPue6Jv08FbAi6zBhT8m339xnpX9cfvRaW+f/rMWEHLQHlwPjzgsA3C7mlzspNNkt1792en
y7/72DYAYcS00c3zP2+7kMSTHCXubEZZdt53GG7D09a6xliJ0mEDqtme7WQVbPWQ4WScHmtG2sKp
y420bsBZWVIDtlObqSPShs0k6F6anhQxywEhc7nRqknj+K5spJhLyPYKd+wjABKqjCRpkNWzwLRi
G5PblCw55ZdH4cRC1zJ5EFtAzcpw+3g/30h35+FJx611/VyIJFPDl9KLZvwv3W2m91qrq1f+M4rd
FSRpXDPmqG38trdRK4XPRSRBDkdkrtxXRUwtGLzaarBYTwnFAcnN6kG9T9/5eBwTVB0i/7igEyrU
J4ElUT7DiEbvfDjHuEjdmYPtxzmLP+1wNaHK33CUoGF/9r691FI2+PAauoK20h/9VrEcM49/m+bF
eJtQEQMU9EDWSiYgwFPdkOSE3A7lOaAFcD4+eVTmDLtP1sXxV0joKWheTYNXy19V5hEwLooBAJMq
W2ZmUYQ2/4eC8fP6APMMI0wgTvyHN+58ld49MJbwUCXDVeHTku75lVXjYToNRIQBEGGZT/VXTY2E
7gHcb7RnJCSDpnohtaE9kYmGPznOJPo38WkWgsvxVGVwFennzk1/W/GcZ0qi5YRl84nnaCY1lIFK
F9YYCjkhw3qVuZU38hPvmzDJUhqmwF/XhdIe4IyGHT+ymZbw1ddzxbPxUOlYYLpilXmYJGT+/XAZ
x+l1NlqS60n51s1Zxc90+z1uRwKU+vgVCtF1M4wZC3rAG70uQZuR16EUUcwdCzN5UZcZQyUrHyH+
CwMUB2bvyWC+RlohjHJXTS/Q9hMDxyE86pvp87XcoQBPC7dUEzqgRuE8Oliu7b6gAg/R2poQrn3G
WQBxyTq5JpszaS2dzXQtx5VYKXd4Ro14qTvX7+Gy2NjWHsbSrU3RJn8tVJiix8ElK5f0XrTgqdhG
l4aJPwRWsKfIaqolJSNUpWO98WV7/UsiBNAp+SM32bTKuz7UeAcpIx9Bx+ryjYc9Mwws4jONusnd
gDBzv9rZsAItsQZkQ3ArRmhCv7rEJOpKhGX0KZ8vdHn/uy4cWMbCMF6PUQ5wV9LRmNiVWV2w+0Dw
TEcGYm2F6ZNcgOGD5yk6Nlsd09PtUSAPXwsNlt4/oDKY5zWR845SrijdO3XMEytCd2M+eafblUfk
StLv39fx5T9P5ulEHntbPWzgBpayCK6sygTc65py9+qwl/qhDxjakABHQpABAyHiNmbwZ7A5CuvT
4ugXLvaCrLoIw+t+74TnS0P2t6Q3bsAE+YhKr+VbEQwoMxac93Pd2XYMQ3/I8tMwjY2kBkt2Bxcf
XdB4gvNNTojYsdLL6Vl+fhx+X0dkQ1uHKF8nN2xYql2id9Sx3pX/1BjgFL1K+23dcAGXegVPgp+C
LIZEq5kCDFs7802WgtO0DPT7t65zAdul3T+IvaaUuRaDBzEYCAg+LsWTEhTBgplLwpxt1l3Mh7qY
YjuSDko1wS2WdN/nfskir9xD2tXB1BFP09u0vEYlzHv27V1ZgFQepHAbOXUUsOK3hAL/B3cOH8Iw
2GhExUVHFZKxbk1NRQpBJpCHJrkANvE6IBkyA3dxX7d6Xp1ZXo0KF5Sdg5Qqwv2ygB1xr1oh2gX7
ill4X9PU8voKXhvK3F7oQj0tdyI78UdsLTzG3CV80y+t5suiLmnkm6PBFn8chHECQLPegqgfm/MX
6ek1neWZWmnTDq5sH4oviQrSRXW7g7rqyUSMrwgjJjLQ8vuXudM01CB8Cy0ZBRXdoDZYeYngE878
Zt8OFRu6MkrdcZFw+67wX6TTPdJFh9jQHPbDtWuYRiVUdJpfkdkN/QVX2KCUfWJjv4kKoM9hRrRQ
KHJXRYlVOL6crHCQWyeTzjDryAa1HemOozyiWiEbpdfaD3f0JdiyqpqKCjglYQFRZMAvAkDOZgsK
wgLBo3XDCzDVqP0Mb/uowFSxyLg4zkNntW4xBqDwJdVrN9OyixrZscWCHr/wuHJs1DUDU7QEzjX8
RGsc4W0iJ3r8BO6vsKw+nK0MmL45mUaygF3JRDRHuDntzHQsObLHfZ0k4HEjWqJYphG6p5XwPwK2
Y0KQEVG+dF/PpDOPZif2i0cw1/XRMOMqKTrH1EWXGB+QltPeYz092IwkOODproMnyfxUF9q7Cg2B
nkpq1AlSDdMHMLIWrDCGGWKl9DGCVGZOko8HlA2SZ3ojz2+DrFEhrys8Ocdjcc623Rgwb4okYfmE
pPDFG6Q588AksZroJn7T73Dsy9neYslAMkI+ANgJcr2VxgarHDLsK1aF45JO5egtyxXLPz0ns/Bw
oZRYwEl02JHMe9XVXs8KviEhB+0GCYAYXuPBo7HhPKIAkg+CKwhXYS2E/X+phiduDEDXGauCFZRC
zmZhPsyDlbtl0odSyy8Gz38fFHWdO1vQ993bHWu6NS5f12pA3Y52WpnSu9hvB46iaMFvL5gytkFv
43sxD4dtRiUjXQq/eLZa4lE+UjYkfcZ6M5S5J9k9Y8cTEEoFhPFR7/vmnLEso2zyYyl9nf/sR17q
4kRbEfy3VKxGdYT2uPz8WepxyjxQD16HefHg4Hab6XGWHaVev2Ehemjy0SHZYc13D88w4eGzuhdM
2CraKBziaQzzaGGq+RwR1flzPOTbR9Ec2KwF0ifgzQIJqvLxowYu1f1U0ygQOG4b/STDqWUnDB28
PsAtRrATieb+n4MLy4mFQM95hN5988Gaw53pqr4A2UWSPwfllTdgmlxW2eYjM/m9+1sQK+ar1HLV
+hpfXT834CALJgldn0p5knhgd1HZY/id0a35XVbODojEUPwk9/by64OwDOcZT1SsoazdqZjODBs1
+UvFkeRuezmtUjCOUa+VsIrkvSK2eQGmcqvdmM6dOadpG/wm+2sHe1Xw3hp1nTmtn2QOTl3nQBRQ
RB9+ggICVQqsqDCjPcocelBIzX9/QiIOyOJSE/DRpgzJV/KE/pmFRR4VEPgNOqhHbmbATwWdRUKW
wOTI3qWIvqIxlVIZFPNV30IIK5vihlGOx42vUDu65znlLKKLK7+6nMQE0jlfMJNT+WogTSSv8eVf
qqAERoyM60oLJ0g10iS92vySLqvaZ0DqZHvt2ausbCMFLi1O27UD7z7IRgqQKAsMiEVNRBKExQcD
exmJOisOcGfT8R+6gVWocpFTKSLHL01rLU1ZuBvu8QmG8rzf8Kvypa+MX00RRmHKdwncdJap4h4b
7fn/Ic1NzXdDXG9ipFUPLu2KVr8yXUJiy/darmxBHCyjnPgyK8k0XoMCCyvYg4i0MJWnq+ywW8tl
AmZONO8+7djWN8E1oEhxYBOgdHfDPbxqA2hrAw4ylpRyZDfLE5lIbJNf9BlF4BZZiOdoy7svpUJK
ddwZthexei3JT1XpW8UOHAw+ExCEB4N0E7zR7FP+bU7WphKF88u8MqPSlyPt8ek6VhdbS4Z7jv+V
KqWlHb9TXxkTR360ltcwVPzvHjewqX/rWMwmGFM2fFoZPiS2h2u+7Y6MPbTE2V+fE1w5KeYoAg+e
U/BSz8xFxlrHkj5vdyXw6plb3qBLbr/VSpt0q8S2N737FL/cfTTSH0XxT27r3S4QHoHZ4zpDLRX2
TGTSsOtgjM/ip/wNuYqeETiowSCcFFTx32CU7nN6TBL+nJ/njWHi2rPgRV2ueSuXbyMqaiYijCLz
Pk0eURXbkK3qqxtNCfNHqZE9LFKfATY20dYmBMHPCpEXPMvAtVMKepgTZ/V9FQiH0rHKVsYuE2bl
Ajq+hFxacSlLrI9QJcfyGrGN2K/IM7J7fK0BWEahb4F+yrVGx265gc+lZaXnzWIOgnfDy6RnncGG
PlFHFhxHdpmRZzLZvFq1jV+04NANHL95W1es5F808mFXBTN11qLDYiEjjkX+KN6GdtFK5QWhPaFC
HTcp7KZ1uumQmmzuBao2RSyOYbNOIK0n9Ti0bFTA6doIqfnTQjCZ7HOf2oq+7CMC94C6CR3WLYkw
6trnrxK3vJL2YoK1sx7oLPI4nM/a9o3ViddQyDILJN53pIMEioqiT/5xR6ECxXLlU6zXurB643N1
JNkVwUSw5F58Is7ZcLcskl9VXFxIvLq+GXHZ/9RwpB7udNBcUK+lSJ6+sxUZi2SX0dYqa4NqNykA
qUQZkA4de64TuRfdiytwx3hEBAeEvUrcKa2+vTXkCHfGBbYXAi0OVvb06Q3XY3kyAXnmhUWWUo2J
Z2Y9bacHeyY2lM2+ggrlXfVK7sXbbkpmMIxmAcLTnHEyxI+4WIY/GOVnPCkKkvngPQ/BnryNKEJR
4l82gxc9tMnqG4thrm9AZ0RgI80hLMQaD2vIxynu7d8WjpfjnTmwGbNE4ejjtRXCn1p9a/Dhsk/r
VmL7J5druRn6XYrMYqjLgxZ5AzRYqgD1yQiHDfaQ01z5qmGzFNi1HxB2qHkLqCB6HKhFyGzfr0WU
2U/uRHWlQIC9x39/6XQwU98CAvf6kcoSwans+FWKFja+XN0fCFcM9yWs9+8FPB1yPhX5yWoDXuWf
eanKFMNkuzmVThcY4oqvFq0ZjmhFloJ9w800AckFwCMIV1rN9j/8xula9UfXbMEXEn8KE3gtDj85
Lg8K4ZfVV30EBl+Us7ZO3X0g8AgUU7RzKGTPlMh4udScEqqyyFKVLoDJNqP7MFLD+B2wT+l63dkI
SfmPU6dkBljU26iZ/rI++9NMOqiYEZohH3n59ORimmwrAPE+TC4DdI1FQ+L9ijtFkhv196JPdwXU
eIIz2FQe7jhSIrUjluw14Dba9snmEVym4n8t4352hDFI5ivhtdxWn4DrhbZuTE4kkMwevaQGjTGQ
h6ihD3KIBYdkB77bSlmNMmnWEMAume8j+KMxshb+wcI5h/eMQBBUApjf+ocOyL3/ThJL60W5/RQp
wlOsIVM56l5yh+Z4PlM91xgwpFsuV0YuFdZQoxR37KV5a1VrsExrUUiIlwJpUFJNvSTXjlvSuV+w
59xXvDJJ4u6ZU5hVq+KH0Oie5ZDx4Ps2CAC22gonloSJ1APFbyUFJUoprCFCuwZwkhzrjGgCbc4F
bzzdWjW5y8DsY8dOIrjvWKD+Sn+zV3kH9pxbJsdbGcX1NciIB5Hv6Cgf/vBRvCyUBQVz62OubGi1
TUp9uP8p5dDRLoh+5JuDrZE5mjNabT1a8PTuz7gXXsuyj2DP61BCOjAcJ/qLZrir0iV0GyGqy12v
I3TPgKXnx5uRV8aJIHVlMJnUhqV4nTjl9mwEhqTqClGiQNI+3rQyQpPeAP1B0TDDktS73RtTlZI6
BmcblOkjwK3Ic9iwXk4VJ6cD/ziuVZxETsNSDRiVQR0hTjkWte0C0fbfvp1aFnknK7ciLooX5oWH
Gi+QVaCmRRU7w4xDeJVrc7hy9w5hXZcdPpMPzMfau7u9awAHpZTcnM7s3hdZpMCZAq9yZ540VZ30
sQq5ahyg/pqfJWvvZf43h5Qh7ouubDBpVdncY+Uz7rCua/yQUjnQaLvGrhO+nJzhFNuz/p2AESks
/Uorug12yYhopKv+jFcZSSuryrs/GMNNUTMdpBP9kaq6oRW0EzjUq8nala8wHCjw879ENN9/MYop
VfQd0Vf4qpLw6RtCZkS0DwhCbDbYrIVK0ih7mT7cJYZi8rqHSkmGoVnv1M1hHC119b0pqBJmea6Y
iitghvvAmxjj3vrH7YZU4LafRaWSO916Y9w0vsxUZgpdQ/0lafXXFV5FqEJvVACLYqrcQXQyc3vy
Kj6Q94jm2rSxPCqiArZyZH9GKcM7lklYktItS9+OobLSke0x9JxfLHRJ54NKQ4YWayqhUwfjYZRL
oGttxlAJgjXusD1MXACSr/QvAoRAEjQ3gz5oK0xxpk1G8py4OibFb/4eoPNS4yqUnJswX/jfsiRn
gt9zkHomr1JRFERoPv3npdD31s73drWCo3YGzzuJnDzDvBwCc26ic+MxEroxGuhfDvr8usmwimBy
nBPI/bKQ9Q8b30MWiTls05klMo5Q9eaHzcCmtfy5S5eaYNYNf0UKxaX2Gyfgta3tdaq95V894APn
dSDTs1FhmX1G4xUyyqLn2i6yA9PwfNfFegvBKzxCPzO3jaYJIgTmbIF1JPNR08kIXphTGWJTWjh6
Z4UcN6E7Q1GHIc8mKP2VU27lH215GBJhHr7Jeo9mkFc1hIga0S3Kv9ppoaCjjt4bVePP6eeK2MIh
9K3qXDzb5HjhuDhmQbAI9qxD3RT21+9JZwHT8kL1Ex7vsJT/HKUE55zzMpPE/VCI/7t8YyeO5jpt
mgMVnFljGxtZbKK4b+jPXv44/ozi8dWpxFNAufW9Lg1nEyuMG2shDjvLD0ZvduMSdx0G+pxE24Hs
luIJoASVLeHm4vj5G1lG+Yd/U8k5vYuly2sFDqEdeG7Sfj6enHWpQtIGrOornz0Y/k3n4KbaFfE1
AEvOury3ZWl/8WY1a3JFykbbFwyyN6jEP5SRbeWOLowEakNkZr2Av2q3P3ngDS4J0PnS1I7MK2zM
ntW8N7kukUZvDjTo0gFTGNlYjRo/ZbhVluS56MbnFEivQS+Dp56GWN2GWiEUpCcjAFmguLh46tZl
ZrRkyBKTmYjj4x2sdaOnD45Nvwq/ois3M79wR1yQpcONo9rH6U9gx/XOYib/D03FHbBL+/M/CRPl
ZtYhHN+ZGiVSyh4lzTIy8hpDYjESLAPwYsnPRlEDNKaRrtLTqB1koFU+1Tw+jkREO1n7G5iD+t6S
EsfV35pr/6zsaC0mSRxaCV7zGl9G8JeEGk/P+Le92sp2Nn9ME8yGmy/195ubQ2G6yXO0fZRCudQd
mDxN55l4eyxJYYmFTGqf0l3HoeEI+pKJjyZHDVnGBcFjm8w8H7vfZ85FkdpxYJMEb4aJ5aP+TiQe
TDY4MK+WAtDtNHzpqlq4Y6ArthKlol7iLpPTlu5pKm/CUVvvwU9+hG+qA2BV2KeIaEBYYuSkq3ds
6ADp8zHWkbMF0yZJH1b8ccdqMn2mxBrHtzI+RZJK9Pym1Eok/W5GCqrA3IkrsIw1d/ceuz3R9WI2
jsv1a/pKi8EHNaOMkztMV5aPQHBa1HqUKf4LLCq5/RRG2najedWysix2n3Q3sRcya0uvm7qjwlNA
IZ9n6qxuGTz0I8QtQKPoScYu+nWVIgUm+EzFzBd2A8ArMlcpLbC4wFlBoM5Ix9sdsuDnru+B2CPq
vlZ1LCq0Z7KDbPFFMl8sdKDuEWSKCjff9xxyKYuERlPinEDpjPoIzdqwr4gcU+tdAdINo5zWAA/G
5NaqoJXtNNp3JJ2FRhFnd3kQhcdlC9eDCnMUJ+stl9AiDp5YCP5QiskpjNxIM01sOUeyW4VndsYu
dXbtOhoGKPoa8CRNfOgGMIIb1CYhF3wVcmk9PmlQWAvGgRXul1ZaW2yezXgV54yKCnu01UUcD7nl
HRiJlQxuSGs6mXtMMXb8KBpe/Kl8MMpkQaZXvnUZJUy15DXuzZprGoZ6DQWklFZDdDYquLbkQcVE
1ZIqmsUTQOHjcF/YYMmN1FjwZFIPPRdqOg6zUSz39JOJJwJ9QtIA1ICX5vlVQYFAn6vhGNem2ksS
NFo0imREEMNTD8MoNcclVgD7WwYVY0cDLYk6lKioPcckBx74XtgPdJWjRJPRNC1ug/4T0e5SsNxb
dNDV5p0Ym7KGz5bDwpCPaLdfn1Umydy1Z8Y9GQycZVe10j4oetPg4nh5FEAXOadL0K9x6rU7b3RZ
13rnl6gLtdpH/fbjjUsLVfksixY1WxtWQmHcSTUADWBmY+MDunqP0Mu18ARw3k13kjNAgx2tYC+A
qIkfHbOa2FfQtZ16NedyBvyd0LOVpAESV4zX4uPzeMTL7WD+GlZ0q/BvYsXwvMjUVVCHRcHjy2xg
ikG0ErGUt3TzR43q/hQZK01NoDskDTTU2Aff4s51faPhSCvOrrSuM5Myit0YLAniAAGkkEr6iuZY
EFlCnEeyghb4emvOeK7ZIfOH9mBz6Jhbjz7fO8g3YbpJ2ZRBbsazUOVYupyrIagyQcyOqeSutx7x
GCVlVrYDbedGkkL4AEh2mSBqa3UnQQbOsGIlHChj/NSxTrTaacVZ8UeaBMLCcjLzGXbcPlhFwDpS
wCouZfDaKp8QT1dL9uPg4fzIYe/1n2oFuNYIArsh19Aougl4gjvvi5Hd4NaS5rmfU6jwxnc1slNK
wlzGNx6pt5pRkNzsoYg8FzhPg7oGr6sDEbWcGrQQuB95m01bQwllhrPn4zUVuFA2mvnrPkdQb1su
1VEdrX0upAEJvgPnATg4tlEEp+SfJaFhVUxFRtcb6gYIQ5YxWld6PRi63FoUhQVymG3TjURbi9sX
6WbxHfPqSKSaA0Tgzl60dMYpHfhfa7qWNvAAqRPy4g9/4r7seCGvhXSXhSmYsZX/jBoTab3VeboO
OFsg+9J7W2Z5/nRcU2ECuiQ1MYCMu8EaST6CK6H56A9T4ZEGMr1BQc5GzzEKXfeqpyBilejitKsO
98mSsN3ZKxb/hFhiPGJYwkRzIO0Z1d3Wu42lQYR0VRY37rVuUeNPCiNCPlD2o4vJ7tk/pjm2pYrZ
Mm22+DM3zBBy2zlpMIqG4Wc7xkMiFUNOM6SdUp+a8+QynHlXnj04lAy3Wy6xqTSvzAzwuYwPwMKW
0b3OAri6gAcMf2xe0hI+2NxaJRe/EtfRzDUtzHQ4VcBCLSG02T6g+Ff6mmi3FKqqqoIKfoAtOuUm
of7Y6ObBiaH3By8J66bBaO3L/Wy1/jSmYOABnImrGqfvQnS+Se8ys0TZ5fdC5YAWw6mgk0TFtnAU
1KCE3nET+C9LygzObPsbsrwEBEFtq0zlfbrHjaTpr9BfTpBkc+9nGgq7WwXPo/2gCZdwnepbMOvR
QN/bXsbItECZWuBofURLDWUIknkRqYFz4gSWb+ZGDKKfuJfOcKIqC545CJD/f2Py9sPAOUptZaSl
SXxqKFczgJ4oFwoyPmilebYBPEGv8Pd7RxVG2j0j1w57ispxx2KHMvhEeL4keKoLrWCZMySfNYtB
NTJqnjyf6aF4cFkxjkaLtQXP8nrtyi+unlrPM2U4dqrDqGdNRCQM9Y29GvGUyubghZw/ZGDE/Zqx
+Jxu9CH3XgIz2mombEMMoK+ahdzpusYzIdWfiIaSXyrbr3duLwFkr4WWXkNmOJhyiUYAzVkB6sG+
eqC/wIFBpowXlfYjATOHiuOgOwoqYM7EkQ3F/ojVBFENDCpZgarX/aHv8BvucZtNLP5KBfyCPn7h
d8teFiH6KOJXPuLckDyr+/unsUZivR/kNr/1rAZF/V6qQfj64YhDu9G+DJ5esQkZcZewmi6z1emA
KZIIBnCetMEBqdfvrooZ/aof8Jlo5ppYSFcGEO0zAVsLD2QWK5Ua8/58J3uCXMEfjHf2aEJuyA8o
giydAktn0eSDO1dRGfLZoN4sUl4Yyd71wIkTziqyXTKjRAupPyRbhNK9/yjcN1CFig5TdBbIbEX5
GhHDwob+MpCNXdTrqdgdppW71YngC8fVAx3l5pGaFummvSmvBC2CZ9b406AoXQo3lj6XLBaVZhNx
J/iYf6455RCGZ5uxCme99rv1jLuAesFj8SyFmgBKep9+5h4NZXvzvFZqZwVw8jSkI/dPn5RjpuY+
7dNTU8ONnq/8WMaHTki1cjviMetamNArHjA9Z+k7IvPgwPIBtw5MyXW3sifmOTgv2eAnfjbVk0Zc
HWZsBXq1++98nHlQgmu5IyewY8jt/W1HNCwwE4RaZESv9iu9kp33Seg1iFyUwGmpOdJ3xxt1Mf+2
/Vh7xkdQzuf4+FqhGM51laYStaF0tUYuCdLeUwsqro2+L05pw5TRXgAms5qoYHgtUQTx2DhRpg3V
cggwSkBMy2mNWlUxSLt6QqnFRSYKi4VgT0Nf1BJvuw3v+0g+4XcuovQmAjdaHQeCuwxY6XAR//1N
V/ZdA8kA7gJ3Bu//zHL2KA5b/ZG+oXKZ4UAuRHwSYZ9Y+/RATQpDCKVX3yrD5i4VgxnWaZgUy9w4
xHKI2BbXk6iFBD405DsufJp0vyp0lLrJkCs4hz+wLysMZnDV2o54cADPC+j8bphrR8bReHkJ3hBa
KsFoJUiHZLjROwdcFY349ebLqS/h0FhBZEt1qc9r5rLmY1EGcMC9/ts3HW7LsNDiuIDd8ZYzdY7S
JvIb4d+q9LYwUj5mz2JBJBqvMmPm9bZRBESCm2GKO/NfXbiJ/dEiEEeInOK/c3EBEqAKw63+fPRg
3yTgDo88cqAvn6KF95IookzAwydPeHQ4wi6V1P7UyysbcbDAWZtpIGhUCHnKlWZYE3gG+imxWO9Z
8qXuDaj104g3bcHeM2z35ZPvYL9XMLAwvow+zD1OOA89Hchs2ztmEz4KeRAQe0jM6KOF514W37nE
Ff5W1OjFvc4QkLeC8KZcYw3PTRsoDNMJoBLqaDXR7LNYIZ7dRVbfV8qEYinK04xr99Jpr4kom2i9
zXbKgHT7kjBQgwclF4b30Mv2hN1XJeOmR4crVQbKyFLcBQ4HhtpMiXivfHQwwRHSKV1Jrm+BvBeJ
t2uWnFdYp+nB1LRuTmCyH34kk4jurO85siZixH45QwWIBmCnUL5pm4MTDOVqY9eyK9oZahB8OJdA
IgCfIa5KsWJSNeIvIFTWK0PPhApHDbbcBr+zI6M/yzwac/94VmTxVG0h8aDTNtl5XuXScPiuUC+p
Di0BZRmAAaigrD1FPC4kPxe/ZlEQ9DrFfsv+SvBLXLkY+pMOer+jXWOIgTYao3UJN9LT5F2v07H8
o98CPDD9gQ5Rk050hZe8PwcW+XNI/bJrCQTvxq+GuHttS8c1D8YsmovqPXfEkNvjaTekc1eRACk7
Ruud5wGGI9b/IyPf7PZggAUL8+90gHhNORs5e4yXcPQS6ccQhOz/L+hyN1wrBGqw7QwGRIcm6Os/
sAX8VJ2x7tEkYT6m/UNtc5lxWe6jYzIfGwOQhu54DcRC3boNT5Z006RSsOwNK6YOMQd/LX4+8zPw
HNlzQRMrNzp4ARV7cvqt6ZFKnKC6c8O2lvBeNkWCji1grILfX5d4ToapCsp74hc5kwxepMniCpO9
MtZ+fbSLP68deTBY0vbYStcuHOLuhrdOrYcladaxp1WOTae+nCRz7osL0gHHpi3lsCkS/PgDxON0
eIf7XgXen8AQMd1ROaoRB/wsUlhDoCaM3cFNW9PfjT3Ix7Kg+G1SmstUuVDdj0M7qMI+ttdv/FwX
fXQgXH1tQWSSSdxxrvS4mziYHaVta8O8hVwNzu8CEcgxbH33c+AoqBKGHeLvwxcJ6AxmqYTON2OQ
bWkYfRyXUdkFa1Y2u0a3mLT02303Wn7QnOQBKJVD8w4OJZhY09Kdj/Yiil2EO7m5lyXFAL9WsaIy
R2pPPawZh4IHSMio6re+h+b4M2x/TcDgKpRKJ50PcN+rwf0aOopSQu72bQn1UMquy83MjDpGhMY2
30NwoFIti47YFY3OSiT85Fc0rQiqSddexjuEknbRpH0ow0YpShXqqFW5/3xiPNYM7HxE8/X5+Tp4
91splR+M9jHLBS14mBzNTXn7hTYz8wA0EK0v/q0Kn8LSz8VoYHko5DLi9H9Yw1cdgXR+KShN/+ym
CjI1s7n00K13NVUoNE6MDatU/mrbsjdkny5uuRtuMwzZW614ZpVnPhk0KjdRqONE4cdWoEPGavK/
blhT4NEmPLA5+cSrY7L7Uzl81OOHPX2Efar3smSwMN8mWt4m+Z4QrJh+aLIsaqIejbo5zWyoW6S1
vLnqyw37pf0bOKgVGdx7y33pbww9kxXJm6kc5ATEbmeIjIesJcgY8XbPD0sd8F7zSE/6pHL7kGuh
Lol6BND38FPltEKJVSzOrE+4gRspiy9eceb0Ijqx6/9xGQ+UxnSDWjLEMHeBkIlp/suex0Nrsuv3
Cadvg2WnptNmMRKGLSgBo7VFrPYct2mSfKasc8tE+iuBpOBhbr241mmMM4izNOVd43JPJe1iTNbq
+y+m7TUVCsjaEddc8fUdgT98BpTCdca6Vwn1MrNri5+TRBJOcoBumvJkbbhA+0K1YGPvaAyHScK7
Zs4nAA3OrwdOK8DLeajq2VjLQRsBZeOHKuGuQ6b5i/1iSoDZR9NJc85uZnw2lGQ+5RQghyjEJ/eH
F+uyBA2EchzpeOaWPsT0SVHL+G+xeL2929oaC5ME7T65qhCJe/mwl8M2orDBP+PbMBcpts1dOJnk
/nnLvvWfFqcYsI+fiJia+m9zj7r6MKPdPCCZlLbC/e4jvjYsLIRIkZ7NEOQJS7FDWhYb3eB635JH
TNqWZ6Wwb3/pjG3pZ9GQ5RwozezzXI6K3/0NW+Ol2abkD0pvhnEFY1Yau/wdwNF44m1Kr89npe2i
Ahb+iuZvMJi0AEvL31CXFSCdF4RSEEaBayO9EueINu7mTtuKMPTNHFWM16rZTi9ztzyMIr/nNtmq
YW3u305N0LET+xEbDfSO9ay47EuHw4oCmeCv/pHfeibhg+QBjxNR2GYvHa+OcNCDnhotAynHC4sP
Xa895ZoE6njJuUCm/C2OZiC6ef4qPCgzFJd8oF61dx7C7Y1L51aWpeL5tz2TImnhAhXfFPZ3xNpm
AZOoxyGE3XYlACyVdHA4ZN8kBvN/LPZqONlTkxTv6WgbvnWKkNBM98GvFWWFY7mgzr0u4uhdinfx
8prUP1l4EDQFswWfnERBY3rNk4zU6dJRykxX3aADm231bYOm8BzRr915F1Hw9VYYlupBBQrUAwKH
wj0c+3yDi5WXKbycuu/JVlWhiBxQZ6BvHD/VIW5jS8Zt/4D6TNrSFcB4EUuVftnTGiZHc9l3BKlw
lDhQs3yQcXIerrc8iWOYK21PIwYF8B8wO8wrPZ87QKGXo6TvFBEsnqDOszVZVJ3mqz1LuqqkAju1
31kxbXCDhyrJ0H7c0IJgeETB0cD3Y/CcB76BWNy7HSKNhZ3QFdVnATS0DEBIiIPiRKKmdLaCKr/y
hrcuGSaLaLLohdUCACBsYX4xd7Z4gp4ig9WhPfRqSmr1wAtZPqvDFtSaolXoyG651fNqoLtfoAu8
hXvg+4INR4kWB6W4lLIb+IjxcHtTIGlnbc84Pab6vCajy5OjXlWWYBdnXg+RhGJdg6mql1yKRVPn
FeYK4EAYdUxgz0ISqGZ5efUU+X+hcfqBt1YFmtenG5tm7dicxIlNhK/q54r3tCNwGeEP7mTKH6f/
TFITVpruPVG+sBdhBIOm6AB+sYgwlxfICmBl1AUFCCeSnLbQgILaHUU+zdW/nSUwsa54KLJNLeSj
AMMu0c3RqugVCqCh6++C9UjmNHSauLG0kXz6py8pSJqMVEbsXMF8u9pE9aMRlIdz6g/hHAH43mE2
e9u4zwSGz9Bp5rS0sko7WEW/eoqqPa5Kt38z1GUz8o67xjYas8oOeOZncm6avwaScrauGVEmCmzW
jBc0VOQ85qEZTyVHjGtHdaSGJkbQ64FSirdk9QpqRj8XOt9egkgPW47NMxCDy5fFUYJ3jxeoVl/8
LWHCYQWI24IBjHTpCuuuWej+0S4v3SLxP+an9/QXfWdQ9QemHWeAfM1e2sHQ9I30u2PODAuYCZ1q
9yOPKktcnR+u3snrURkmCwSs8Hd48pQZyc2P2zLJpM8fA9/Gms5upfSpyQ4rmKgPgsmCV7Y+Le1j
LyLtkuslmPlDDGum5PhpyGpQ5BmsNhPG2WV4gqcxQKAkdfuWCyNDsGlG3oDURUC0Yjq2mgtjvcsG
Lcw91yWdD26YSGPYbx9nsif1jCyOS09yw2HjrAPWzKP35XIJWAmqXUNkP2DKZIfI/U07BkPAKr89
1zdbYobVB6hDMRJDBe7c1nX4cC51oYVIbJELneEa3T1Gb+cnXUXY/PvTw3nBW+8Old9jRM1IbI/J
HuyO8ojphvw43gA4o6+DpjicM1Ln4J7BfWzS0szLMvYSiI0a9koWEvtYk79AVTXJzHONZaHgbhds
VvNyeXoy0MVXliImpEdcrq2B7q021XD7FraN6OvZ7F3sR7+hP7tQunRX2PSx5Wj/4lff5UpbQyyL
6UHYY6rShOdITPCcO4wg71jh+V6UYW+jwcRPzGKKjfa67Lx3oGD92DevQTTsSIkwhLxsD56zBKCo
iuN/WFKqcbbUoH4XqTwAMlJzx9HHAxEnurw3OZw4XB8ddiquTCzg3hHHKEqHUVNGwUyD7DrrEbn2
0JXJ6eKbmSqYaNCU1EJ39HVhyJ/QSKy/JsYE2gEFqioK20ZgBI61s4y2dLi/SzCJgcZDtLXuH3UP
mmuADy9XAkODD7D/wXFp/W27KHSJ8KSmEm52tgg3QGyL5Fb/6apkCb9GijMVF+6KW10mokkUinT+
txBrsXlMs3Uwv+iOOqyiefl6XTm0XXQQfwTBZHLMxZpwIhAZnFhGSJluP6R+3nTno9sYU8+mWZ6Q
0WJMqvt/tf4I31zBbCX7ru7sH/o8CIBzVakiuq7SFwYSt+tIszPhbCMv5+R2cBdc9DKFOr+TIhsn
55cv705riGKOj4lCdFdqwB1jqBVtdI7jpCd6+15YsdGF5l6aWmLs968pV5h5iWcS/Lr7eI8zU56Q
RiEbgYY+qahe9rn9LyoohV8ewH3K578bCq2tqY/INdG8UJN6wZf1EGpX00qj/RSuR/ermKlURLyb
+Z9KXUg0meKCjDzGBPErjmyAxLXBBHYgwM/tKC9zm54vaDns+WJ+/twDNUosxVwxykJONKcAvIpj
FyLbRHA3mW99E98RsNXCfnLzbSVu74WbnAfjcbFKaKKOKgWs4p226iFJ7eqwgw08GWP9CojIjksV
9XW3n+Onxrx6zA+IoGxj9Edjey8Y1XV9F4yXcJnRJRjz6gs0Ek9oIKxhq1kNMG1xQ3lOZlavlrVV
ZzAG/Hs5+SJfat9AQA9lWk61yglMjzUGVCDz737F3IiNkzfmAB0Yccbso0NwPPAVPuMxwtik5Wpi
Q9zU/T3ETZcdv9FyRilZ4hLFlCxXfKTYwHkNMFXySra4UYO2N/kMeJGWB3d+ynvLb3DTjUiuyMRT
N66Eg7cHZUSvOghmOLZuIbLSpUwszdfqgnd1+mx1JlT6xhAMnbo+bfpTlT0sFj/hyxZyiYlCd4zg
BFbt8ZKwuA/ubwwwx3uMWMbgOSpOH4eXgq/VA1HcvLdcvBL+ZLnkHvETJVe0O+u+aRDSRCRehc3h
v6p30ILt1aCaH7BecclVx6Gpfs0XAYbJmrEbwpRrjFh4qJbVj0SjBCU18OCJJCL7NBg/ehhqWfnC
Eck1AKutnBuTc815COPDJoplEjtQkJSl2U6S9UHRbhCS4lQATi2442Uu8rGeIFa4C+2OZJzkCZP7
ZDjgW3oC8PaCATY36nE2ybH/ZJF1yYSCzS8a4i6+jwZMa80FxDY9uGsyqPZ2ncpS+YCGUQ4vWdel
2O3BmuPuEA2e263ftraAneb9H0l2CcfvS6VwjIvGtYlb2f0E6oqNF80j9/3vXVqt68t7m1C5fMck
kNthpBqTj9fBDIEUFiqEG9HhY2uoyz6huN8qwVCTUvUHossEzw1oVkcJQFg1uBto2JNf/1uCsqwH
i+tA7sSfl6ry2cMCgL/q30hJxTmpCZXEoKP5THemAwavKkPuGyp2M0dubV4GqoWVJe+T3aYYZ7Nl
OQqqUVtCgikTnT62W2/0IqOqlwruo5H6e0edPi07aLGMoRzANN41AUOH4DMgsrUpP+fEde80P4nX
3gt0W6P8rONgT1Th2eBMuuL8PtM/0KCTb23OCnVzXzBU3fcDE2xcGUfgGUsFE75OS2Ojq4yJWPna
RjmUyqO7d5J0/+Or0v0hpLYfFUUf+3FyJPzKCOzjCA2AiJ1jOBvRpDLcTwDcLhYLYpQm4U/ir5xL
owvNpiGwtXq3+yqGVulRCEivj8PpzrxFmERwRW+38dRL2f7H7EMkq1aRa/RPOLfoyNcTgztwkzzw
y6bGGwMuY8k1iZ4X6/wSY/qRjedlil+XVu2NUPaW9HM/3tgyio6VG0n9HGg6QmlFSXxWC/iaXeLy
rn1WgmHz5PuTNfvriSl+Kh3oLQ0BRpJDMakicYPn+8fXw6TElTmGEprxgukpKz5qF/8TWBQ4GvhL
4iLS01y/BoEw0ZvkWisonA/LFj1ZXtdPnoaC4GUR21fq+F7S1CbohdHfR8ht/9itO07ZSDAyeEmY
eZ3E5JC4z+9RjvBO2lVOndEymROjWMVFVJwgTzsVuL1/+pNCOd5iXaOlLlWyr7zF4v3mlJehWFgH
+7TumoYOxIQulyV+BjAwgVXlh3YGNG2BQB/PGBCNCLgtH5TuHvagfBojlvdPod+IVEDpRqfrvPUg
flY1FOn9Wdg5ZTTFcAPJAnw0lc/pOCzzTCcA++srYKPlkHH8mbkz+dttcuyzBJRckar4Yd6diZoo
HUDa/xodPNK32cbtx3LySzS+ldenKr7/BXIf2baeVCr9XzPHxN/H+RmqjJtsQNqT+WKvDqnRG3rO
ghqlCC68PwcjbAIy2hVMCXp0nN8iQuDizBCJERwdUKz+8Fg553z1Xw5vjrijQmghLjbRTerHOTQD
drUU8QU6/o+uwhTovonlDnhtNYtxqpMbNV7JK5E+SJBSUWHcNcsOErHESNJOcSp3Tzer5crdiKzN
NgyRaFY8rM5DI3MQH/BVI368A4DqIb0yH2vUmkxtHm+lFyOibxPcEkup4BWRGWFcz7kQfD9OGWwj
z3cB7QQpf5nIPG/cfIeJsPfwnTfbR0JWSjwSEcB004TH5vO/dO+QXBn1IwstjVzy78LG/ZMqOfJy
qtAXPNe2ejkITDMegfGXhBuidUIWB1EBMQcCWQLar4rg+EpVO0OJmYGxvB5rBvyFsH40U6b08tpc
n5+9O80kpxQF0lK3DbDqLRF2x5hgVnPHxKpWqIiN+lprs1XhBtMQTazfX2C3I9Qab17+KLftlEEf
uOnV35lFbtk8J4zZ4Ncesg9furN1QnRQ5OGzobKYyiLNPG6D4CRcLeOtAATka+q/9zaiOfkSW7FL
lxvUKA/BCFHO9Nc5LCKDdb7uwE2Qi23yiS3U0mo1v75TBp7FCGj+aum4AlqhIkU9hYKCacfef7BD
2bXFO4/lwauJNgYkR+1uZTTeQPs2Fl6c+yfC/G5rbfr2kKzVj7+/vgR6PYjN9ratudLSHIqaUbsD
Hb1EyNsK49TusatPhjdvD31f9ggvokjzQsMTamW+wFpx+FtbqWsvTb5d8wZEG1hI4MeAg7+fKrul
+hpU3gC5NnBKBDEMwoQY9zse6/ADezawVNUjeAIxR9MdCqojIPIRZV+01p6svxiJpvmGB3ZxGWyv
k8pFxdhwI2yT+Mj1fFASTsPg5ApJfwfLBSfDs4rAm8pSbNOTaSu3JF+wWBu9h5ghPG6c3k3LlsMt
sMJwRgKIy8E6DngwoSdoKb1I8y7oYn4mGwKbsqqQBokj65rDHl/csob+mejeuty2EOsXpra95okU
jPstBvP5Qme+/GFI+qYZxKJmvRzwcZbiJepVLPD/BoBv18NVgAjxpOQUH69R197ybI19TksyUifp
AuDVuPwAFY+IwwhJZhiHSUWXiLunMcEx+3d+xr5ggohjdM+7bAH5limWH+d/IL0Hs4BYt4DXjWUb
hVooX9foPTV103TlTM9/VO43hO3FMYWiYIbOGvSFW6thA4w+jKGdhzHcxlhihRQJy9lM8p6tpCfK
5DigED94jqgqI9aBJvpZpc6WWRiMeSe9xbOfMjjSa2JLOjR3VQ+2n6vbJYvsYX6fV61wrj8BCWuh
OiGaReHvlIgIBJFnAAVCUW1zs/s+s94MN054Go6pqWEAOzr0xHFDCAcx544WIbxr+H26iGDwVEVf
CEezcJy4t52thyFWZvj3isowCFIQ7M9X8qUa2O1k2xpb/3Y4SIIxFYWAtPbiFHwH0EgHYtxeRBcL
s4ZYb1a9vwk58viSyU1JDVU81rizY5Ief4z4W47FnN8eNu5mDAUeenNrH1NhrMWbylwIJQt9idRV
fxUrMQiS/7gp0GKP/MywjZj+p5MYw56gvc7Mx0t/GUB4Z7+rq78BFfw/Ul04bqcqiPExM+o1hX3W
THpzT1JKA+pkuRsxZmmuv/0bC+5dawJ2Q4RydSQ8Igh7mwN/oTSl8XAbBYMuuoZ2/Qx0w80chxX4
ouQw0JmEshePD3Pp7C5cvgPxeSz5TU5rbP0PDU3F053kUS8Xd6pVfTjtTMAlap0lfGZS9aO5ZyXQ
FPS6e21/Y+dUPX8LAXMS7WaASW8WPY2YrIwOEmFD3ruJKo7kuQdePvosefaZyuAB2yu1mB8SaSwc
b0ja3WG6iSgd05fCzOevI6nL3VK5ZiZz8RduGIJkNuPZ6x7yNEz/dkDxh25588fFAZzdFpsCmiHI
DWhGCGL+Wi+Lr5SgVKD+jOhw5OkfBGXSPbEH9S7IcxCAS+Unvq2cTMOOfnqOZx3PxhAVbKGHmgfB
TQIFe7d+oFZ/RfwqIPeKm+9tbLBQpXJvoVskt+eoPvkilDNX6KWllFD8fgHwvQJ9dKpAKakBmpp1
iyA3teuk1/SzxID5V0Bdg/3oIuntGWWPtz0s5dGrKxtYlV6omzXHwulFWdPeEnETyqKIzDi8EwUY
5A9PldfJzSJHTJNOjzPjRCQRWeqABn5bI2vwi6uQWrK4ybWHPug4Jba9vNf0783a6ED3hF3SaWdo
oz3Ia1QtLXD0T4AfpRVgPQWPaeLdBdffWBDZ5LruP03Jh13/NNP5iKSR4xXZ3wlkpjrVVF/17q/b
vqdQ2ASaJL/iIlET2YLRcP+cp5e4UVl9lQ83E215erWaatE5ypn1wQfM5kUJHw30IT3uHpVgIKBE
qsDPglF8GimyX/DS/8hc/wYfRxluaVQeuAXdKBAL4YCJLKfCns3a7fjKc+l1lj7NN4M4GcB+RdST
f5suOPVQtOjiP5anbkb/Mblx3U5AzugWVxEIAcN1nsSFLC/2VyMPKBUKJdK80UYp8lxu66CbN604
HXIhB4p7RcPh/FqE/IaVpTK0nHsjeMLwoSFE6T6wrcMOajCexYBWqXJVGTUxyp7EpzHJDbPVpexg
pvAkE8DbZJicYB6XI0EtwvQYexGQhImdLhdis+Njgi8UgzO5963nFDxkW6IxMoQbjxftitlJdhbY
cnDvvMlQPA1FEVB14WZ/JR1EH9mTpzHvA8jGOUEKMaMcLPU5JGR+5wR/OTPbO4gzfxXCRbMRyADW
vQO7juRF4keO8JL+vBhZqtYoRsmm5rhEjmblBR4DAjpeivZHnq5kdA5rE4ao03BBxxnX9ZngAwtr
13bqmVP5Yyw9VifR9B3ApoV9aD/TyRJNT51rRq6RDul2xEFr2lhxnjak5v1b5MNFTK9WESLRJenQ
lapB08tlKDXk8d/QuJkDBj3utzdhDX6muKlMidBEO+/74To5SirxrvJYoV3dgUimHMX4jQ/sUImx
hrrKeS6wkValWmuiHc4ov+6nFUjeCWjXLyz+b660mhlHsLQoU4PTqAL6IcGKBU37lBahOMjzTHl8
4MlUm0+6LN4ClNA2kEvMzBT3QTusoKjVMPZWAubM1KdyIJmN5pAJdzvf5KxoFDYiGfOzE4FN7wmg
M7VJobsnym0Yn+/VPFAJVGtmn5dYbNAUAaaTrAVh66hS5oyZBaYKPR0VSP6cP8sQZYewCwzY1eS+
8haR2zsH5ShWk22qbvW/YIvQX9AM/fMaxZNJ40H9W42mjknu/JGj1RnwC+1Uvua8U0GxE8TJLmsS
1V3AdK+iD5tjMA3qAujEZUcvHTOdav6b/y331hm82mwO3ubUnrO+6L65oElSxr3QlFZfrs1hCTBf
iI1Hi3H3WUq/eYrhKSPYiy76sFGpvVXt9m6RpDZymJKM9C0gkgNeP/9AVRAt7T3mhfP20HdZMY7y
XnrqzExIuXDrKnea62c1xFmOj8dxR2H0ys6kD3thCJ7h2UKI/LOLegGD7EKksTxWY6sA+rz3rpBf
Mn829BADLRREjf8/LJUmx/RSL7DdE1PL6ZTxCVmwGWJKuK9XpIdSYZhDOw7S6ZfEuCwI4s4U1Q9c
wE8ldIYPbJD5bAdES31IF+SG9xgXNLjaavtxKNTD+1J8qX69dYz1AKYIjJr13THUVTdVSge6Zphn
15YFvqf/UwT0q+ipnnpHE87GWWeV8q2Pzer0TDWiXZW3+u06k8EKf74CDfowNJLNPIx/FhdjNFe0
RoR9+LN7ZIp/Bu8WtX0e1cz8gyD0eKrpmETFt4Iddby+Mq0pY3SMHG/Ye4G9mxrJQTbdmimU9V+b
HcZssB5PYfo2wxbF97VB9rds8/ce55+3w/cBAajUjwMY5XGv2Q+34ZA9VBoS0eXrFbxMegXpBTui
YgDblRZXc3sy/T39mF/mH0BbIEDmkkXOdYjvE+aYgfYzF4ogRCDnw56KDbS3vxckUmk1k2XM/emD
WmSn1zokPTVLcViZXOTil28dAhHFY1jux/G7/LATwtbxOnv7L+2Vr+DBb2DRmA29yjpoZvpFYCtA
Y3EjaYtDrrfAeBaVIdARooksGiRB1wCVEt6at9nIvvZhTonPf6uiARFG+kC5HV8vcyiw3YqY/J0p
KXuNWLHpyP2CaI6ozrq8IVF2yPYGKudqEggbFZ7rgzGzPKV9qKh7BvbHyc6vHLtN9K/JFw6CFDpE
vDTtod9/NY3L7dFSD3PqkVAH3fqSRslrAz2/dSD/ZKndMGhTjVfmQ7FEdhQliSizrcPmNIpXTo/z
rm+fH5dvHkOmYNTum1aojI7hURmo8XBzs7diqF6K8wbmacsL8IpEV9HjUjlEz2TvVG2nEZPLeSlV
f9FRZ5RI2yiBHE/zVO7yy655G9iwi2ipQiFjq6NJ6DPZnxiS+uB1DpLFnMmJNVR65Vy3HMZU8xBF
9QK0RT8wnjJJ8JvpqmxhSYbNEKVTBYv5jLxYPSEZfM2hoL85GmPfWWjc5Hj++chdIfcXhmnKRMcq
2hHZZfOV1bu6rA4dR47VItII4Y/Xx6kJSmGXbnFfSqEIpsLkiKgpwxCUTmDVsDHYhV71Vkrf1DIT
X3DKVPRutv5EBBn/6L9D5gIFfHPEb/6/bNo4bPx1ERgwX2WoSILzakprW04mr4Z5dmjUn2RLs3L1
9xEm3581Xx5QYSo0z/VlgrhI3IBL1L1IIne+JrFdAhcsBOWlYQQGcV7fgRanaupuGVvRgOYXERaA
yASmdHA6YE8qoacg6QUS86SCefoCZt7bttHIP06UhnBmqEDwpkEsRzhBcjBIzBcLLutUSOEGuX2c
yfAxkFpYF7KwKmGnJZj34xEeFKKV88Yvf/7GKk5U2ih1IZU48Bf8F+L8XsWvjjVpjIJUaA41Qn9X
tibTHAcX3R1NrruqPPT1JhkjEebKU/men57onAjBC9Jel6HxQ8DxqcBwp330YUAifsvDAJlU7zgr
9ruse/+W6Oef4XoAin/LnM+hG8opttBOMEL+FGKoljaSj6vpbWeogijryMi4QmUOKRKQcTua6xmY
+DQ7qA7m3EhSA54XzV1dwe62A2ckEHBFi8ZLSym8UVZGxVJepJXHn+SC9zH+Yh3l9WPB2TJUTI8U
88ubqW+RVZ6OoxNurWDUoQ54/PU39yZlklz/h/NKxosvPGx3XO0On0tOtSiF60dUK8OvRQqRwvh1
O+jKfCO7NHUrnRxQI+o95SHLpKvB6M/5RVhIMek443fLw/cBalAPeYoeopqO7JVnaX6HdS8TURHq
Wo/6Pow3tjvBU6pCGuf151NZbQkIykz5oSMpkoTTwQZQfGNgnbGzV3ae8OA47rzQ+gVFebI5ogoW
mceLzdmNAf0m4HJWN8e/1K8Eq1awmLjAD4EkqaTIrYSE7RBNzMj9I9DeuEvOsjQt9XDcrljuj+p4
zh1uSMGd1Y1JgjNeb/8Y2F6QT0+Xzse6jbBRP4tKDar6jNfh8SEPi+oVkMw1pWg81HSsFf6WIgFe
4sHLZpaGc4Qizk0z+/A+ZqljaYj5e674gUt/lUULFyR4eO/1S0JycyyktB7wV+LPJ6EKM9DHwi3w
LHISlcwbx0bjYFjndRe+vh53kKOVvJgYdmHh/u2o+vloaH7+Cs1ZQ558/hqQz53Ex8G3jmM57JeQ
HxXFRFEzazPcQpGRoQ7Y+raOLMzXu+5Sh0Bb04vsryPfWI9qXM4ObrZ8+of8Poqcs5g+NR1l+KP7
hbJwZil6qeINHwc+nTvnkyv26rDulNH1MZmtZ/TwhahP0B6Tf1ZS+rdYO2g9mn6phUah0SN4lDSV
Hs/VPs38opnJ57hPuTT6kKVFwOMoHKMu438kVwjeCLqxrmLYuUAi0MmUeJV5oqEffs+wCCbrKX7J
1z6BZdehH0N9CjQ2jzZ+pZHxZNn+0iEG8uDLh4I08ALHe5nOdog+Y/CHJkvllwmWPWRTtxr2IcSE
TLUQvUq2f+QY1ajIt5kmLTAfbNQpjBAIyciIzRKadYqwhFVnKfR4YMmdmaBIndl9mo8hWuNbugf5
tTbADRmXatTkuNKTtVqMt140+2ESisG+MORkcVNwll/OIagzgynHBBP8jgQieGo+O7S4cBWsgHfI
Sjuj9Lxq+yR3IFgC0VBIRbS0rwmVDKTbne/ney2Wm+xorxudmthEyNWFq6hSoDeRpSjMaV+4pZKh
6ZeujHgYR3gfitXLedsGuiPYn12yxrXstaEjAIM89MqNZTLiSmvLpvWWzXoJlooaXbG7roIOpz2K
nTcrOi1n5K0E4mLcn1kta1obQg3zPXVmhsxKISvbeBR95RIDU7VBMNg0ci+k6gMbzkKoylZs25Ea
hZdHkyHaGy6wgJr0I8ispFOyTy5RDNHHLC8m9qYcFhphPIaRj9JiWNJ+ARbZTvkPJpKpJqaEuEjd
AmcmXNxI9N8kgFaWC7h0QO0LXye0yDkzuj9bey16dwHekOIamyn4m0VgLR69JvIYocVMTTOeFkgO
PyIq0aVaNAleO/wwAny7A//UDRj0ZpksoN2q5nRQ76uCKAXPNOaPvZ4lsTOHKYg3MU7WOLW5n+d7
36hkID6y2xFZqJTppjP0oWGyXwc6RsQKgzjbL5gWMaayti7+WYPsgvPv+WgZCFOFVqFbmX9bIYcZ
67I67BbSpBwduIcCmmf7KqZZFPvuiOxJjirMfqQIyZjVqOSPMIIq9z25LaiIVNm0AZ8fYDoQbE6N
gLl4fQ5vxEtEDKS5jMTaB0KmEh97EkPf4qh9WAj6NcYo0XkIhCoSoyidm3YbnYFw/101qbT5bVnE
7y6eeB+/PlWSFzTLLgyLqZM8iOU2Ey1s+GlhGZ9973sCpcuHyuANUYdv+HzT+zGTicx8Z51nsPye
rY6om2D9KGxWU6c7Vu4b5lhpNnuTpRSQ0U126AtQ2xX/tYA3tiIJHMrjJvDam/zgSd+EFTAfFqOo
gp7Wdfljeh6XoysGgJPzsHQriyA6LqS+IefIpzXf02lJimJRZ16AjpGdsF9TrThoESxw4vOYqfcD
FGWi/jgbmULPK21GgIkWc181SMR9ja70eoB8j2T81xDKUI0fYlvsfAMcWNEkWhZEpgbInq19DArt
e8tCxX4tySEFiI3JJtuavW5JJSLtOiWMPPfMy4fjFWOXy3a4pfxjty+lnisJd8Pwk2gCcvxhktKW
9WLTllH/NMNhYTSLzNVjndOpYH4ObMjBvhr6pPdX+thLODVpxSimMsXP+JZEX1Q1PdPVV8rJCNFp
9p1gP1W94UqAFUPZ6nX7RFHomzjRyhNfzSX8zhOzzZ5WtzAm6NIyFV668Ek94hZsgnD3GGepsKdm
JvLESRY2pyPZ7miM6vc6Bju/KPzSE/ajodmPKcqzGIxS7GJr3iYUfKLbx2hm+I+U9u71MRtYwnNJ
w31MCJcI6A0HzbNurv5pAxJ6Gs3bYp/rloo84HccnyMYzH4889US9/xfHOmae6a38jggtm1qDQ2s
9HjwYUKdI8EX53+qB1U085Al/BTP19tba2fAN5qnmUCtOGgW8ZA6nCGUvuWErpeUX20uMuIG1TK0
6X2ggXNTLSSWmhXpIhxnN7R70i7njb5BfhnAxBD/1PeW6EYGnpTPM2BcK1Sdy/aRb7RlOD68pgJX
a8/TZip7ehHliV2xjkuNCK9LckxM5n7Wb4JZlD97mjZgU30IpGQvoAtWIFnyPktkrvY7J1Ifcn6a
L3Uu5AeFev8/Fq21RdaifzytEAVpcxeqs9u3/mFgjn3zROC74qIMUKNxSaGFJNKV3zkHiOTeXnN/
AWcRfHw0yUr2k7XpKyp1ibsgRiCg3KFUsQBGwCMEzF6O+he17flVNm7akXnBB20zQO0otg6+5+ry
pyxeqrdShQwv4nsVBXhZhuxOuQmtL8EUItJAkeRlINyrvkI1vCrO77etezmNDJ/sNdgmuyoSriuG
a+x+H77Eoogn8lt3Jt0MMx0HPQY5H6k/WW30jBCl+xFJSRpo/shdKj6lXUb11hPjCLHRQl0SHL8K
c1L35Cr0eXGEPDMrgpwJIC5fKt155bc94WtymXmAOwNvP2vTQPOzYJ7cC2SbtayS7wLLipODghay
VBbSSOb2ELNLplONpbQzyNN25m0vxKkzigYBCD3L4kZl5DcJswAVRTPxsH41Bb8OV3EOOR2HClMr
cToczQ6uRwRZ+2n3qhV6ekXk/CEY5sNtd9ht7wntyopsnZacZz5lKv4tEmPKEsJQv7tUHbw4DVwb
t7QbioC+YhJ7nPWGDQ9IBT4/9QCMi4mOe+aGthuThBm3saAdZxtVvmVj091LOeJs371blTXn3F8g
e7EwLi+XIIONQdKT+LuA0jTlFEcWMikHuL7+NqE0hGuE8Lbj9HP44hlIxsrndTWb+F2XTahKDOIX
0n9KaulQ/dbbCDYKalWGYCoRkvvgUqzfmAYp4/rSbMyd5MHdfqaIUd5yQ0nck6OcV1UzHW/ue7i7
8BypHzEL6wuCY6WJ93fkj29pMIYbAzGB8oQTeqye2YkKFX8qh8wvSbPvZhTh86cOPLjz/vv6IvF8
yIgf3hJRKiKgceEDpQVxAn5rkCwwRlbo+jah12pRGUuJON+ACEXDp7DNkx3vghYdDtKvt/G5rr7h
Z9qVTRO3bF6Xq0VMvZjypHUmlPQHIMF+IPd0Y4Dqe7PiGxwMn4i7cf5w9ZZNsyN/4T6ExFs8BX+Y
i8hDrvh1az3b9/orf5RfAfh0l2vcJKL5I7SZs+GW5CdytoQCeBvVE5Gsn0jDQUh3Y6/rW/mLBuCq
bxre2s83NoauBLWjzw0PygmjQRX44OlMbWLmrIdKczbB/7qFPruhJqsZSiyp82viGm6xCv3+y4Dl
KMAxSVvB36IfcUAQN8Sd6OgfttaBWOa8VfqitfT4FcBldcXcsP1NWNpCjQJGcKbgVwaOlnFaCD+Z
gWbhzLlXMUNYQPn7r3a/NeBMCzk84sZe+yv2b2rDUtVUrv22h57RrZhPmkW47YopPsHamdGH/VLB
AUGKe0d9sPpgdn4o2F+sWdf2SQhtM3LUGoQxSGYDcjWT/i2jdjHvthpPMIBFrChL39j9K8XL63UN
gaKwgv5/rHZNIEnvKP3fVBaWJ96PPN7te/aYlE7gJn2/uWCMcBZUMXEzPL35hvqyNIljs1iVXbo1
R3n5qFb+MRT/FDeToPn9PnuapWZQxp8Y4jD+zilI0wq79z36wHRxmp1k9Pa5q6/8c/ziahDg26Tj
cEQaTr/ry2oP2ctNvZVCklVwEiIxcavAmlSikWg6x0LLw9KZ1k/05aGwIxa3f13iwQrDhsknOKKW
7/bNW+StiRRlr4zWRIlG+ef3mDbFNeTt+J9lYmPe74af3M/invdv/avgsgmlNcj5OiuQc6oqjsKT
LrDu6q5t9st7on7ZQhIxW/DyheVDISh/TYa+I3SJgmD307dgPzah5Y0xg5XmwQjGQ5Tl0scCR/AS
nFLM1OGw17nPajOHCZiWOTaj+2Yu1WT0dPHX8/qX0j1LhaDhn1Qo+rnyA/fnGJx5pv1cyKgQMnrG
CjMqf7aW3h8yPZ7NahyS3LGQqHsnvHAA8+M6KRstE6y5z36Wnr83TlKUr6GPtgMP2l1Hcwmj7sBh
Ffj4U1NnaUSEpJ4ym2KLfWqerQsl+uXDO2KPoIA5ILZwTPBdc1C9yMlLQ6OPURag8SQVIiAu9Y/I
34lP3pzqm7WVkIorsStEWZssKMFssHuLifxBW8W/9dCaXcGV2vE4seGnfKx0ay5qTrIleZdcZL9V
/2FFPXWHU3KbDBU5gpbH+liHN7kmyPPvqILL9O2SmWtUr3GGhiQSJK6TSL6SouvrhAHx60HAk6wA
rdU/vLQgfUMJxVI0jq5f9XonZNHaQf7TQGZb/I9EXPIDHBdVz2Qy4iWlSL3CHxm4dzyLgkO9tNQW
w6HuDHvLMTciZ4KvVy4JeZu8fOY+wz+ApBQrhDGTqE5+bIm2iTO3RW0d+KEOPTSxMqzgg7GUvPCf
Vay3lyiafbO3OwkBczif9tNU68bV5gw5fU8gKyBLJMf/RvLI/2MEJrkrT9UAmqmSuRGcRQXGLUaE
sEV7nwnASyif+2eS2H8J+rMNrKuz2+aPr7e7na5RfazNobdKtmZBdnZFMLJ3jsICLiIURE5yTYcu
OKNQumkDP6aYc1CCrNyHa2GREeHjM+yGwfcX62pY0wcp2zY/bAfyDvON43AFBMOCWDOO4RG7hRGb
0Rp1runouScBUV7/6eZN7DwrnXRNByLhd6+bbjtDGGpbKhqeYnR8qpPS40Bt2tjupo2IpzHulcoX
pbGnjFG/0XkQx+JtqWaG/l7zANiz5RAATiDXVZLM6YOLjMZFBOvvf3PfPR0LifD88ssSyWbHPA/2
UZn+6EJ3+KFfrSb43HLeMI0RmW91pTsGuXV+6kQa6WKuajEiLiivLyg4HmPQ27Va9AhL6LlwkY3q
MJUumucX17uVsviMJR/0If9BPCzh05Ab/rcG8oDDRsgh0t6+fsb2EHh8SiSj7b2cVanAWj3D7Wzb
xOKBM70w+TUVxnywNWDo0/oS7788fAlCS0gvqOwZcea7jYWwxx+uj93dUK64ceKZ+rHmBC1HP/4t
BBCvIQUzAd88Mtxs1UxcWOHxBl74tto+FBWhYh6Mue322HhzGhi7dw3Oqnh9ubCvBj9+1StDEJs+
O+mFed+hBqRtQu2/k5/wGiPqJ1E03Bzrl/BkPyLlGVVEISkIlEKftKIFVHzopCMKTE6J4Vro/5dF
QIRUKpACkqekLRgLjbni/2+fXxz6n3Gcrbix0PbvXdX4LZVSBF8kJeNbfV0CA7A2T8Qdcc0w0sng
Wak/S/oyUC1fWzOQtYa3DyLIxm3Q7shUWwzNaaWABK8vjmhprJ0XPkVb1cLesBOjEYXlosPFGx6l
1C2U7rHQ5EFnVj/Saxrl/at171Jaj9tvnnFmiv1AAMuteovC38tuRJOqMmHZ0dnQulcsC5U/B7uI
ZxfHcC3hoYp0TQTdVd2UsTzqcZwLyYiPPZXBxqoMm0KsqcWkVVmp8m41UuMfRyOyCABoMbkNggvX
LcyRZh9VtJR5MVxEr5aMvjJ3Ktwdp98wUb9Mqvt10XlZGNkYn49KbFN4F+yZAXENgxbzLkrhqQCJ
Jt4zAWBCS0/vHstlzm/6EYfSyP9iZD1mlE2Eve5E2lU1Sq5FKBnLIt45xnxq+HHeSH36xMOBvLfi
ietOVba28bsYKbF/H060GAtyisHZlREjlzEElfGVSnRv+tdwla5wKZUnoMNKUWCMh7pnjT1tlkyD
JhhLRwm5vXdkYo93EB+5yzGz1Qml30tRqu77UW0GXntnYwtM68DbdDzmyoBWbslcoS9juN5UWqpM
+f5hLMSdBOd52gQCoX36+FhEcvIY4dvOKFr1I7IU6dCuMj88HiITM7DnVw98/Gha1F1D50BTb8uD
HvpZ28s0qOyHOnvZRCWn4pGu8e8Ufv6zMXNvXk2Nfrnduhod5mHfzBpql8XHv/xOH05Lv+yS0RhV
VX5LX/coqvBx3ELRpsgWNIGpokYzs9K0wIKXYMZwgFVH1P494FQpd6XSDtGDgLV4exoSWhhYMyAh
SPMbkgzAsmRlLmBkuJtPySCu6Vyr42t3NEE2bmJZE/ZQkiQFSRPzf2te2aVFr995sfedJPe6NRFR
edr721m1lELA9v487kuuwOCV5f5OhhBuQsrXgm49vfhIbPoNMfxdva+WPQv9A9SFYNFeYgHX5638
aHrUlWqwTMc/PTIzBscvE1aeIFnsYYbhDOteeKGjJPqXRocX//xswwJaU6QvNtSpXK/1oAvmBpTt
t0AOMVDwY+Q+n7H70KiDTxokEXZ5mKQq7GkvTzFXoV7CswWKKbHqcqlfU8InLc9dqvTH3UddaWEa
HsL7QEQ2+n324oYhKJ+cC4FJn7p4QnhhNoXzVE0E/NF/YWHRVeE3GMdD+PyMp0bGScwHDDKZ4LQw
IUfI/RAENWsuLDxtQYwbTJj9mhiaiNp4c1MKzM1M9KDBYbQHqlFfMv1dhtlmIc5ecIia2Qf+4SB1
3GOmBvcq9oWrsjBfKLV71j0bTNCXNowTrfxcmpA/08AUI5m7lhU7G3+jkbDXQiBsuYTEHqfcpnlD
T/V1krdtKIDvCy6u2rzl/Eb8spzFGc5KqNH7jNMHh0KhVr4Rh0AFpZR4wQ/tzqKeo+17Rlq/6gTi
8IGVk4vi4n7BTQcTG0eApGmtODwY0KBTgyqBApMXCFUfC0A85Fo6f1qYluJWHwj3Sy21N2DN+pkM
qE0gxTwC8nSbXBctPzSdIO6c6vS+i/W4hPN1WEPd38dJtNklFoFYap8a7XvfTFy+WfLx3evSB0yJ
8uUfmSYbhOxE8Ve4Jiqxdi+X1gytyWZQ/nNnj1UiB3QlbeAvmMX9dbRYGugIG4U7a0ysYtt5ClfD
ghHvyQEHfrHbafQ4aE30D0RYMMqpShW2Lrq0Mpj8Ubg6S3QKe059unyjt4S6LHXouK1Vf4CgtfId
nCSU1gyukTCg+BGVSOpsw6f26xDq3w8AMCYrXfzjLsWDRWaJu2I4KCfOCsz4D98SjchOxQXYTXud
y0oAH4qKkhq6jzcq6zIt15g18tqbT6TLtWYBiInb3bWL5/bq3xyX1v+B+IqHIJ7wxRHOAU9N7T9K
GO5gp/ezhmwykJpCATQT38JQVw2oFp06akbTpHf1Hzq+enrh45D9OOlZF2WyQRWtAbN6SZJFFCt8
HNwL57bc/rBj8O12aUxa90AW+3QxAfHXQfpoHavYRYGkllS46H5A8qe3p+BvxgRwDB353y4MTbe3
CZUAhukiLK4E5ZIK0LQk9mV6J9g5QzB/b/W/mlYmMDbTtXwgHxo6tWARFTEw/gMPPKxAF6oKkNNQ
bFipD+B8rrfw8nLDPEtZxx8WlJ4sMfJ1Ry97HN8GAwj7NBRgQEvYvfsocHlb8p7l5tIdKQk19g7L
u5zVeRCsutGr/w0KOLoEd3UMCVhnYGYffehi72wfEF3maALPevlAFM00GRp+q2vYdGuTQdSkxIca
TU6AFRvt1XxYjXanHYLzzSr+CstQUx4pJ0AThBmYfqjvC8TygVjYprLp18DlhjZ8jM5a7FvKOYd+
VQg4CxrZtZjN6EvyXet2CkCQsaVHVXo+He0eloJBzgkQsErbZh9iksavpTyPXkZySYP8gDUgavi9
ikjQanDPAy8Mij3t6osXi/yc7fmo3ShJfzVnrtotokNCbVXkEZkCDQvuAJFEC/x+F+aj1Axzw8o/
FSoDXSDzmLff6TjcdwR4sfBGTA0z2U6jLq2/hR9CoXeY4mBMfKRv3mbtHaGLRcOndg/iyQ2rR4fc
T/i0uMlVT4r93su2X8skxUZGKVp1z1QiEL8fuxyGoF/re8BNwJ4Oph8bOLe4AOrfgSYPA74nA0dj
31jN/YQQXBLccBKe+uotnUoMwEpiGOB8GESD9WuuVXQrhW7rLtClXncqRYpFMkm/ep++ra9XQQDe
ts5ulxLk6P+AoP8dTOmitYVRh0g5+WS1QIPWHr7ioMj5qrjnnlMxezYzKWsEBEl0WnWVqwQEIjOD
9clChUAbNiCQVSW/++tFzmHI+b1vntQW2bP43z9DzzlKOkxe1rPS6pNkOy8d575q8R5BuDTN4r5i
7dUIUN4QSCw3SmtUejVFOrSnXj8OfpAskHenFfmtLuPqh2IYETLVLIiwc2Ax5YL4DLosXAs03cSG
BnytWJugofRml3chguljGFob17WcpMO3ACwYfLklP2fZ9eOAw4SIb3eOG9eFe4tHKDDaRI1GAJbh
6Hz8AqrCMTUVjl6hOZKNRhWS9b5j/j6vXWyyacOOmmRgmxo3Rm3/4nWugeBejSq7MOVdE/D+FVrI
Hp32iA/8+cP+jxSze4xx/+XtF+I5mHCOUQh9QbXwFSb2RKbVXaSySDd3ABJqULOVrjGJAmgm1Ska
vs89DKzV/liZEdhF6afFZjVcRpAt9Zrehev3tA/RbEIOvdDqZwc8fB0lOzyYVMUB2pjWBOn8SPZ6
EwJFZuKYGO9lfXd2LjYKbaAPt9TnZ6lk3PpPYT78iH+XG8k23AnhdrPERP293Tsgmrw9sd1UsAw7
a4HhX38l6ehhm7ph+EoBZB7L4pPjBz5sK8d5wu+bItFUIVIkZbpGbpFZ/cfbOmmvn5VRFUbVPk7r
jNY7/wr9gXzyC6RmAKx2npr2kvXoWxr1OIO2HLI5/DNgffS3vmYCcWJGCrj8/xJWNyLmsYyoYZ+N
H3NWfBSagSHyqvQTTFWTp/UQQprevnePv3yRTApfLMRdZTiZWJfXoc9Mj+n5SkJDgOfQf0wP2Lbh
e0R/Ws21Ror7Ofll6FVzRMTUhLwr5SztfhEbn2YqO8YZT/1MGD+pIVgGMBI+seSyD5xPob4NukjG
WEqRMVLWj2cKIx4LlHKodmD6O9UMyDprNd7TrzyyhCZZm9Xbys40jVx9HG12puodczI3Nl6z4QAE
+9ou4VEUo3tb7izYfdEFMLo/YG7j4hFpRDYaEZaaUnkIZ/njlykaBE856Ykvo88mKhWX/5uCp1br
DwNjj7RqSZf8hpno3icnMZbtI+EgaH8DToE6WzOYhv2H98BzVdN7AKYNODUOkc2J5+UEcHQ2kBcG
SUSFMDo16VAmIcz4yl8Jj2/Z3wvGnucNGTokXaJxngT0k3ALXHEhzXAR3/Mi5MYZfhfoYx+RPLHr
PkeXc9PWlnX8AC+LP8DwxVBUAGTllpPwrXdVnUaXYOl8V9Tag/rRolIKqminKS9g4jolsW3oJRaJ
RG7ulBNQX0d5Kx5hRq5rIkeCnoeljLX4RnuKUpk7Hl8MQvDVqbvoiZBvEN0iMgQNKes/Q8ho9Klu
uFTG1MVFF8Bw7RaankUrgKjRYzO8Rjmt0xn+5KPuwSdSek+olnfkv/zOgVZAzG2qX+Egqu06Br8x
BTUtBdHnKQj9JsTZLQRmsZNmdOZjySHu2Lk6r2JZDY2mRdBJMZ7vJgYBGIZ+XgAPCsIrTSYu7b5i
6QzleZ1S+c69bRyHxYp7t5LyQc1TCzmTaylyWVEz6C+hK9QQskYcLg28MEA9nT61ES8ZwBeXA18T
P41sm4+jv+KDP3V/qafXXMqMuhHw1SG2VeepQP6UlLQlMEuI2AVQixP16Rf6tmbXTic7QloX0EOr
NwzQwSWsGEU44S/j7n6wRaRQoxkYIRkt2ZfECVTCuirHA4rwAMFa3V0XplsgIMzUf1C7ulr24jwE
ctQlR0GEa29KPUjSxn3a4wvnSnfnJHN5w66j7LzZbqDQ6wCBmiH2R97v0t8wOPpc0OsqYLvrSzXL
Yt1hHQWoPzkX1KU20nUvlBZnggloHIob8DqE6pNq/yyx5t9HP+6LvI0xeM70agLWnqsoG4B3KTmc
EJkWgFnzPpU2jv7lAaoiMgOXzooxxAbiMAIGM0s+ZRbxWQIaOI1gdwmL0FHIuKDLSJLAsVh7/Bq9
Re5iZ9hBEt1FwmNcol4XexD036OLkDmdnncaiEteJzASJhQTRigQA16EHYgBAl2c1BRbA954b6ne
HTHaKHnMwErja2qoz3MGXhEBcdHrV+2opBVzCg4fC4VNjaGIDr7eCWUSBwlUtxC9Rnfqhqru1gyA
Snl9d3ri9kKyVZzeK3lHEgYIgJ6y/x3f39ILAuxcN9muY2+vixitM+1zR/Dc8Gd2dplox2my4tX+
VAXmqGDuhD0fWRzTVBKpkY1WuGcZo5ycM4l1FPkRFd07H2z2EIJ+K4hneSNVMXquqimm1BmEM3xa
0HSU5n7Z2ieolb34PVjHk7oVCPSOCGTkIoPRLvl+XXrHn05skgMT11yG5LuN4ptf4/JYS9f5Bd1M
wsE1MpDSL39HB/T7U7jnpbJV31/e1Q3OR+E2vOmIIkX7AZCXy47sJOZACXGYOgEJOgRx8nEwWu/4
u29CopLK6DnID5e3J9Z2nZyF+a+GnJdNkwdR3AdOwrHA7q9b5UiI62uyRs7iSd3W6NpiV0bq0qse
eTF4qKn0UHvm/RFnBIt17kIliDyO8LBPWcfmlm6gbWPI2wenP5WSI5mrQ8TMzHDdGvNdKkOQGC4c
xduwJ4EZwZn5j9Ee/u9Y3Qkofg3XefZlmjcW2rFAoawrE70g4p4vIwyMae2mKJG7yEDvg9B5k3M/
zmHyRYMdgXKyjTnfTFD7gkLwcfGQYMv/hlgloIsYdnXsXMlrbIrN7aSX0cLh+s7tj/GDKiZluljP
TkraU/6mXg9y3QFoLM35HFcroSgCynekfIHg0nbVp0NQL1e7rIDR3J8lVf7TEXVOqkNChuaAEWIP
A1lUNNvUePadHDAh4G6sXpvoxRSuLKNw9oKjXcBVWpzDR9is9+8LslGYr5O5BaqRIQNPx36G0eq7
8UcgamrzvPxyfKnPatow3o7g699v3XxlkmxIFrAmXpChXDTwiJ4bWMaClPeAOCG3Htf4/TRBLycn
cLefd+9IY+v6sb7jYrpFE16tU0Tk6k0jLNnqmLSSAyOMv90cg5ZQ/EYiAj3snffTDbgO7/yKoibm
EBt+4mJWif8d1dApoRqGGwvXgDDlXsAF7/daCbNWS/EEUzIV+PJkc6/Akb1v+bpdp1eBknV7OBCA
16vSk0DeAv4BKaqdWxjlR/GFREolAsaaXdqqXfyjekfZQUcix1tBbgcD3BcK+OVOLQB6OG0/zA0p
VYZFQCxiAllrWekMv4XFQ668KHNyzUP7RG4qyFxqR+W+qIjMIlXgfQ8sp1AF36et0HhiAy644IbO
adqVe/eQ+pcLUSEXX9yJd5+Myy45G2Dw/59V2u8PHUFeQyi08JxP75JIAmSE5G5/KTH7OxRV3HvN
FUi79wkK5C2GlgwLWYDbQNyJ2Oxx1f3BNkOOE1EXyXdsuNT2Vprw3OHPzNEJrPEtBhHrCp36Fdt7
relwr677NUOeWPQHM/pAwwgPWkz2jOSqtS3mFFCPLkuQ5aHWK2ZRbxkUinuqDAcc2WHeHbJDHn5z
H1JFyLQXeT6L9ObJJ003MV74vYFLfOkyAGfwf1IaWkdJhNlrwpHig48TRIlwSmlP6Yb3ik9QcjgS
GejIfwAdtyFP/Q4UM0/MevPnhxVPp6oTKR3yEe5o0Qxhg9OSQ5FGFoiMwMDX7u7a2hYFRvYyAqQs
GQQLZ1Gjk4YHmeul0JcKjUgiz1XC5A/zktWAxHROoh1Tz4AloUHsbX+zhsjkkkvb0yXKg6LHNAsd
0CCCWMxNyQ84qualv2ZDj++0I2Hhr6eyb/qWIUIxoJHbECipvw1Vg0QfafKm3QGsA3WHdwSrm5dr
eJQFzd5jrwrQmDzSrmq6kTNn7MjHWych/cCdw2gLVW8ZHbYx2fhqbJpYAAetzgs0lE3oNbP1Hwc4
hJVbzh+J5p5kcSmKvM+zuDGD5w1ZZhnER5cfl9w//9A5F9nmkJevqb/JyY9syppoR3kdHvHv+SJY
3TilSgjl5rxHuQ5DfMzSnaXRnesEkaC2JgA+2Ar+JbtfIQ7jNj4K4pJ4/7VdQHmF5MKlZnO7wUIr
8RGPzkBMjNpJllKwDv+FRuImFtMyfnuWHWl82fV4GE6o/p8R4jQDP6jjotIky4rkZ3cpPY27/Oo4
A231UsYVnGPTi+KIx0H8lYzrJrBOK/bMKJv/7Ut8b2U6o1TMDFkoWkNJNHIVJHUh7YkyD+/2osfY
62VnhwJmX8QoOeaQySrF+lAHBYrX68pXwJioaqofaTj2UOZz97i4EEfVvgYNYUrF8QABkyMvDzI5
MeTJ6zcNUYsideio+E7XKSCEt2j2YtJD9asn+yedtIhsbtYJQF3kY32Cm0rQXnbF3U6p9UAsy8TX
iuj+UD3m7jGk0NjRQETAX99NoVgDZ+aiYMRqtxbh3n0eVbR1wQO5cvZtLBE3AgdiNLTnMz3tjlXa
JnY+saJfVg4Lvnqs94Ha+ltxJl0PZbMmuMqAwsjp5GFruCeF2CGBTe9ug6Lw9lnRJe/1Gc7Tkd72
aNUvgFCyrA9uDGroq4P9JqWw2qxffShnBNLun7nboeDQda5g5Gna/4SB7cPp4Ggrpdi59atTIrHQ
a41NsKkD6dasuvLTwWG4q5pDoIjKiGB9UQTscPChgGxToSBi6CxrZB7gaH+bbvHD2IdrojgwLi9M
0TNkwt9DbRRdN0MySUPPHbr2g1D6wHMKPZEETgoht3OLpHmiJIsNUNzaf7/FF2Tthpy/ZwRYNPcK
fxZ0L+tN+pJoFi0/MN1/NGWGKwbLPhLcV2uaeFaig0hI3qc7JwDMlcPquDWAKLSSecyfkDn7aEyO
OJDP7/dgHkSiWV/PgEybb+DQOAZY51tS8oAQY+GhY/Oi1ZgGu14WePK6j+r8du8JJWUmoVLz1gVj
AkE3/3nyIwQ7gzAf0D0aBYhrX3YqDN0/F42wKx8HrBhHOyKP4BEaEqGuaUcIFuXuUcrlQrDlGEIe
VErOt6iEWMused6FAf9doJCVOhrNoDv1x27bX4qeY+W7qJC95p+EB+paV3f9bqQmw3yyiGqpkZ28
gShGunSFD+LWpMXMJgFCu9fvhUEjMJ0QBX3KxVw/7DD+5+uyLGrOYtQFEZ2BsPvNrs+RASdVkwcO
fQRLUV8T8+hAq1b7w8IWx/LbMpFF8aeAFSP2lcu6YyR8il3x1bBxy6s2USeA+3pjg1+8DmvCw0q7
rzVWy1GNC6EuyCbG9Yi8wZ1B2b2TiPGhFMR4CXbi+JODK8BOD+PdZK6+rGVDztOuBfhmQ67DoEEO
mjQALB0J5klEc9oSw3FFFOLmxwqiBUZmt2Fjzi29/CyhHYTTsto87tVLuHHMRYzMd9Upv40bXsEY
ya5WBAGqN1r3RBeCvLpJT05B4D/dtCHO8TfrrAdyxL/Psj5DQfTac7Fu4yHyNweGmLrq01Yq0Grc
zDJ8GSBK2PeYnr2n5isi1u0s397yVwOLNsEUoR+NZygTnr14YkGSseX4J8KGM93fkqZDZ9H2TJJd
Q+Y23KnqllfgSBp5cnSguxiJD8t7Chsw2OSHoq8fN0QKIgsZMKS8mY4b/xFOqQuAFaeFwJJtRYxM
S5rIBKiz5UDWDdZA41ndrK87KBuckBbl5X4FSz0wPrlWsPdhe54ZtYSEBipUnFZ9fhAj/Zseyvc/
l9Xmg1iUO7OOclRtD+kUlPethwJjZ8ksBnApNaBy9EGCkWdjJ7mCwrLECp9uuqPcQXi8bfRrAGL3
Mm7W/QancFvXP+bDFkOP0k3Cq2CVoLW4+hHiOQsS4ONJ+94grzOi1KQiBySwUUa/9OuA6U1SHzpO
D6gvD0PEEoFDQKB1rW6/64DDoOe+B2IZ56rio3wA70/27/ayZc4OmC3INDmsotbqKn0HPjijMODj
OxcZ79ehmnUAJuODtT4CsT/mRk5lrIZSjsp8KBTMfCzjTKEnSMmiNjYyRCX7A4t3t+LKI3y1YZo3
+0IvsxxSis7vlO0omd/KL4JNmh6MLr63wbkAYsmOt/k0dcZOdYYzkvzwMPaqr8E8yxTkI0HA3aYZ
WHhmPECdw0L6NUNYYtWIhS4zVFs6qhgx8J7OyB2HMDbhlhLq9aXZZ6LdN27BxC8it9VxFBNBychO
cbkg0K62s9wXRBNzHsBxuUPqVUWm6HEQsELI2ZUfhXr1TDK5h0Ztp3aHoawaREFsb8w4NtT6eMkl
3iJpL2PSAZ2DmeoRH8Mkxz9xxswXx2N4SqXi8+7TiiV48QqW208ThPHr8dfPpcQYx6NIaXln/JtJ
rMGsKhgcNEkLFKrU8U7ltaZlbm/I3j3x2ok9Thip/evZiy4IlMPSEdRzDHB7Dv0aV2Naa80JX9ri
C949HJQoujMnXTVEjr9Z9e6CDP8ELCz093qR+j3jw/I2VTeM8DTgqDAfTgsoBTs9uv1MdKLW7tyx
/xJSD9VJUASRaj5Q/4Y3lxWZUQgz6ywCn4KjolurRaNsy2i6QbIYE1mZlHCXvGlYqTnlyzMKJuhm
0NlKhkI1hi5h+aX7IiJRPcArj31D4MwMcznzWUjSAUe3O821Sxf/Cv4VWSb7ZJmjKamoeSMRK5iJ
jLOK+82e2RMFsQe2M/IbPTt0irbxqM24Wci1JeDIU6vshbIbRr9ofG+AkyOy1TOpiWzlJrT4lg6a
s8vWoGudRfvaSeE1mKLBIPj4aYFTsHBQb4BP8yJ5ixDEbhwEL2dVC+9C2qucioJHiNnnev3aj9Gb
drFdPnSXer/AquY4PqKB/yKXmI6wTIzHpGwh9e5RRp5+1zq3RUHmmldjyrUSJy9rDVDsWavUOo6x
dGC4TpuzeZGQsLXyBFeRKnALvSHrigwMSSGkwfLrtDg0JC/VXDKhF2+KpE8CzGxmv+EIviu3fL+W
ITyYAkeX9YSCkZqDlE9Fhw5sq7oxMpuqiHmzPS13L7acLrsXRePYOmBYZbHbOwsANBOh1MQYFz37
gDSM2KcATIigrL7hzwFE6UrQ0maUdonkRhEDEBUFsa4LPgDvsWaX4WpfR7zyEckHMHJXMh3PCScD
9r0GB00jwOOjVI2kI4sdf/OCkyx9TPUOE2OPuax9p/ZiJwEwKhqlbRQ9UPYjBNa4l2pgzfTkG4uM
uy8Mc41c79pVzhTfbdwve1M/UOq48t6NK3HmXCC1ZfT2DL2ahEkZlUAA9KiV1wVhNMbIDc6HcSk5
LEmME5sDB5tMTQZ/i1CJuIpYEkgVpWlj6PA/6r/8jdcut9k2p/uYDOIoVnxj8ZTzIWUGjRPgwkj1
QMT9yBusjUZL5+ARp6W/04bNuTaJxbRIeqp64xFYSOrvEv2iLly3zWY02p5VdTlP8FemFtAAQDkR
n60pn67M7LtEY89DcwOP/CNkFYTe9M2AZ6E7FR9+SmZe690//vBSG+GZdWjUaqKWDz0fa2bYepGp
ppufN1Xu1wSE6iI4KfNALp2hOm/t9Uw90Ia0/sl/4QMjBeBDSU/TBkYbTkgjPK2G+diI3EZ6a2mZ
jO0jJGzoE0SYeHBmnB8CpJZW2+JQqwTaYkMrqcaXXveBAgueP0Q7ZfrxMH4c7q3cth2uBW78QNQG
amXksT2m+ZxDi38w7ZPgzxAAN79du8Jqtvp/jO0sYq+9uLX/QRKk+Vep2Wgb2WRMC1uU6qIVyB2J
cNMaSL8ViIjfgGTGxY8waok8c7xz6xfx3eAqpPsZ8NPpnvpFmHYe/xn0CdA1Krdl18Rb0338EWxc
2MTYd3BnnqKFy24Tgcy2HAwq4Uf+n5FjSlwkffRCcxLjUd0lOBhSI1NxjdYLxhbQx3+BL8Ouen+p
GPTJdtqu1UUX1aycNTQSVrITjRwu5/6SJn89rjUkkWRanlCND7H6cb5pdn0IWsGUXLUa0nqBoePs
GgAGnTOJtQysyOXL2K5A2fHSYBZ8QcFKDiI3s9+nGmVEdxGCzQqYjX2ZmNvKInednPV+uIhAaIkv
IQWOSwW7mDlDkumSXJJJYdRopS43IZpvL0IMRWlmb9KgeKxUl2+bFQDVbgFf8pFQFqEcnc3FNbWF
zXHJIEK18tsCRnQ5GSsF6K48cMPP8/YM67vCEMYuVV3FKMT+YEqOQM0rNcSAeyF3seSBGmROgpJZ
R+rw/OyVZISVaLfQSnGZB4mc39jeEKlwIgbqiRATRB7VtB3BQVwbSAjR5PE8QQ4/wZNAyuKGd10r
1zawHNtqiiCTyfpbtvDgh3+NsonY/lm+7LWN0E7GtZE+d4d/PZp+dyvyOR7FgtSIA2auyPDdYnfU
J7yn5RS6GDOaRZaRVv5X2vBZA5RgVABW117qDkffHnan62EGyuXxMT0sNB+q0I38H7HS8vzSY3bj
f3Xfxc9uSBKf1pTFP9wVdq6WeypFHlWliTS3K8n+8lHrkh5M6Vck3YSKPFQ6PJP/raI/z9dkqevn
WJ0KaiCSSUuxGH0Yn8Wnrof/EKbMxyToEHuoCZN87OSqhnZa6onWS1R3sQOm4l7sjjbjoBgVcN9/
xJauKhKkAifNzfXjm/QG1Mu7ShcI7D/dLrZPE4zZ4rARj0v+Loo97ASzKdK+YCe+vn05tpHEPCZN
7LW8i8DC+jYkLbnMVgqkdnTn2K679+CP0XQLDGsf9rK4de+ZhaPyzmAKLSLiDAS/Wp7sFdido9Rz
Z7OOjUc49mySs0gTQE4QxlBfo6X5PaQORUqQGUzTsKmNtSKKJfwrvHmlVe1ixxcREo1yZOyViu+5
LVDDEChCCarwTPXDaFqfjbyz0Cg7jlTNmM900VR70b+mzadMp4B5YrOT7UYNTiRwaOmK1chXihjf
7hsGHPwJhy2YI+t/T9mT0L6ANRi+nAcNOMxZUeQjr/sM0P2ekPFy8cZud8XIVtrBW2WEdspvPHBP
r78tKdNag+e7bEDW479DbDZFBeME7+4sC6qLbBOWYJWMYptknTTsLSEyBGHM5hxhhJ/Q2OBVIjsp
lF6DMkdTHFhhF64LRXEc2VfS37OTBVb9pMTi7dXXSXjnSReQ9ZGgdj6LiLKSD0HwfSyLc4U6HHfY
DXSdXiCkEdzx9xKrDDBPi9t3Vl8R2/KdU42sWFKsJv7Ooka5aenL03z+ABit5YR9emhpFC41fgcu
fN1/vMhsMfuyEDg1JFiaXKYTT2FNA3SIrFaOq/CLWwTk//JQL97FD1CKk84WORelcC2kwHQO4Htb
JdbelrVVTE8QEVSXkPltvTKLnpKu8aJUktJTu+vucBj99Xwk35XqofYf0ugalR3IoVdCMWorxD6f
1DC3xBmnzHWhCYrlBLLmmZJ0IiFMOC8WreDpD0qXgJcIJA+Nxfy4vmlUMxsFMCAguA/Pj+8eQ5/+
yvN+MRxT2k464w3uHW2GZ2pjbeqqYvFgsY49GqWP3BhgDJJZ1YdKWfeod2prKjnEmiuFbyqTicc+
hq0K3Jv/KT2UngixKy67bcxnEvobOb9/T1EvX7V+z2xuDKVQSKWsf+X72uLBcDsc6XAVgKM8xRxK
El999CbJz8l8Ixjq06e56n1A5Kw8Kd5zXgeRLLQlKmNS97Qc+zBZT4yvJbss3qAdTBcTVdUPNCdW
V7Okzfc6/S9uf0CVZCyENC+0MQ/8CbV+uOrYHom17IfXK4nM+BFlK10Pd0eZWhrVyUQxL8SPTGaE
//1Me0M1DUPgxwOXaGs42oSfXFM1y4nwShDFHUuOXrtP68A6KN5ZVk2KU/DhwuyJ+88GNMHjjo+r
AQPj5H0XY+p76trzEJ7BjGAYqk6AP8Y0MhXZ+VTqHYLByFuYLClXnD10XjV15+YyEKyl3HlDPC9A
V2RBbDsCX9gxgnuDDwCkoB0OdyJt3FslI5WOje2AvEqkCRkCXkcRo5WTquhq8qT5kr69oz3qz51p
6HrJAVzyPOfrnsafLrjd5H989bOEvWsblVIao5AA43er0kw7evvYS9G/4tOAQbayfsB79Wr3JMnY
mqNKHGVVKqy0m4c0EP1X95HEluQskGIgZ1EjLyCtGvDpvBTZS5iqDVWdsAN+NkmtAOJRy/cI/jeo
Hr38yj2GcCnGOkZ/GJzUO2OT8fHAPtgczgifubGrEmXIv0QZJx6Q3ELPTgBpr+vpqfWdEDgQjjVy
+Iglw7V6VguoQSlv7+s615Yb8ZWWsMTIWadUZWtJXl29V3Av/mW6JnZhuRwz68J1E/e3NnQ++tci
HN0+CeFZCSQquxSb7VgxFnk6UOYc6jeKnRCW/861HUy+xw5OnYvRjtnZb7cmVHVxGAM12+L7TqM1
IW/aLz1gt5ji7GDoWE9eij/gb6qVkmJrBFtT34Xq0UI1+P5SiBvOm89qMvrJAAZrIs6l7c+w2QB7
SvWRgZgpgIerLuxQLoSLw/WcgiSxwdM45WoGzAANP5FpwsF4gUVrKWOxf/QiNB5cP+XvAjhN/Pdf
A7Um/bpg8UKf4NJZFRnX1nmauXc8Y6Zw4FwzGU0cA/hkIg5HJHUV7Yjun3GdQxm4u2T2GMfQ+1A6
xdC8si3u3/fFQ3v0IKklw3q7QnxQcMFl/USlZeYpS0o8AJqeZ2vhTfQYO/KUs0MqplDDwZbFG5lm
KO5w/EWnWK3Qm+vxz3R55/YbV3bburPaWrFEn4fV8kQLPgZi7u8NddEqs5owelFnvJf2prCUlnX6
4f6k3toyVyAWjK/PxO+34hceSYM+IQ4Sm6hd1Zf79JIiAyPhKj3vjkQN4/PVDOctOxGC73D8M2Vg
zU68YuaW/n7BdyTn5Xt5k8CB4zq1Na0HKfkCTF7SBujUzPOFB1h2R82lesJvBaoTMJUVEuaNHrWF
hy1L5WPsp5UAj2RA8pYxAzIyk3CmbIlezutEnjOIvE1b9Bs2YMH26k326jssv24RUjPihU5rE1E5
Kci+DNA0a135QgpGuzufzOPEUCg4HIQK5I9aj9bFRKYD5aY3ch8bX4Ez5M/a9yftC/13CSNNqvsy
GqmjZE7DpLPBpOpd8s1pLMx660b1WnkwD+tpfZvSblDIDa7qCIuuM8M5Qh+7qlpQN0p8nlPZv5Fv
0B7tvnL+PUS0YfcK1Zqjx80L863ApmHRRHw9/PjCzPckX9KQorRVodAes8L3ZoUqKC3ZfJSsA2BX
WiqShXy6NtdX3y4/S+O/i6RnKgwix2nw9sKV6hrUFUWVJ0r1ytVFMiIcMJcEoHmHEF6sxpR0MlgO
gBJCmnTANt01ymUxXW5jtdRJzD7hm9vD7TsoX5eKoCgnIG+iN6F3Lp54RVjKAXOEiqPz5hhBlJ/a
m9NdX5UnQD+6Kq50R6NFAXkXqqbUn0NpL9Wa0u3jSuafg4sfQthEu6ZDc79TAs9E0Vq5QllYAAxX
dsD7zXpkeqsrMt55KssVbCOl/D0b4M81LkVfjONGw3qYj+LkQyD9p1IL+wvC238UDbVO1Ovytd5Z
RKfSrPZBlbD3lOcCb92cUj+zcTTRsxcJSIRbO6vTXpXs7H34ctkY2uhd+xliXZAmxMiOXmAHogIZ
/D1pYIObX15CwYjEYQMLOXwkyRG+g0XUpB5GKhfUrjX5ZalMqIzX/JAmonfNwjJZFA6WznIaLLDZ
WfYVRsw+TSHF/MO88KFqJB5nUPfOmTUd/qQIfynJkXqTHrD8CnPGkjmZngULxGCfeyDvuSN4XXOq
eedX1hoUNcEpTkpYtPPskKcbJzUTuH3KUIMBrAClVNBEEOqSJrjhnh06Mmp+2Xeu55XTYH+Xi3Fc
vHHsY+aWh1QATNpixC2hqKNicloU4n4XAIkrP7HAW2tY3mmUYj68R5GTKsZdW0HUiuDRa93d9Rsa
4drZMFNUjemn3LttkwqRvGHYVpGPA1/1ronVyiCNq0ObmCJd7zM+p3lqtwXA12T69AGlMZGNMnMk
UOjGAAIGgpCPrCfmPRb7fw5XB7GAIoDnrNyYq1D3hSszxzVenwikWW3lGXrXGuJ0oQlD0z8s3cfE
/9TklLMncMRjju5W4YkYAHGw0AMvW0pWIbq39I20nwoAFnNfEsdB4/25pPTBxJo3dcxREtHz2y0K
QEoGvvgU20cMR/bksHSNbWHTQ6iwIfnOxSZXO2+RLChg2b/w6j7g3LJLDqC3SRVdvK8GVtMSecK2
8b7vygnp0Lj/vcQJgs6h629q2p59qVDTz09/Gdj6hELZ4pVPEHgWnRFpQrE29OK2wb3Y4MFxhXLk
mq9bALxO5dTv8TVLxvdehLzzfEDUJ2d/uoell/Q1OtlQbKb3ZdnOC3FVgeOgC/PkZNWUuqqTfrrg
xU5YpqhK5aWKn6L0ApClKSV9l2QII/QwNdPTehDOPLRL/+jdCTudgDzPab3x/2ZVmxDnfMYyFFLT
4tDU4F9B5SevIlqJzvVu0Mfk9Lqp5hDB4/cmhWuyRcb/5Btoz6JbqFURRqqZHAk3r0WBKvOeNGJI
2d2MgS7YBwZIdx9qd+v4EJ3hrwFQKRaku7Wja4uMGsT8X+8zJyH4l5b5cOMvGJ1CtIaXGuNE2o0Q
JZaRQA0lxML2B+jW9TeHYx0h7emntu7yijhxLWr45o4xqwRE412QteGu2jp/DTiB8TIN7VrC92na
rM1yh9SxWtijYxa4D6kw7R8iLKcspslknORUbtCAJtVsoweMzNR7zxEa8M0PW703gXjCeAi7yJS+
01zM/o13S/90+GIJKQHKa5ahuM0IDyhOpWOszo3wuJYF1nr3jVY04l7A5VU5wO3js25KbVm3GQ23
/zYZMI4HsRvduKw3mztHqIPnDnVihhUOrR/wvl5MqUQjTwzskfGBZ6Y1N66+qyOKhivkffYVPwu5
xwH8DFlUFVjBGSAmSdoQUF+2jJ7zNsUebsQrbvjeIXITemo3KU5xFU7STKT5fc21jKrsOdcRamoY
s+0iwrKitixF9BbPuzDzJbjZDZx3MYY5K8+98tVnzlPIR33PyDJm3qf20CTJvG0krgkfc/j8sKG9
0ypi/y/Wu6fGMQe5UiY5z+ynoig/4FEsWgqfStS4VlysArPdKLx1AXHQUxYUDTqwIw2dbrkBcppj
VZGXmQrlgwAd6cvkyZvTujRQ22FZwpXOKL0JIPrnl/sflRiMNZMcH1sD1onOgutPnaxvsckQ1jMr
d0u4hvfGtcDbx7tl5wbgBYVCtgLx5BankSvgQED+8x7WDtwufZgkImt19Uj1aCRU4ltKnx7Hme+9
4XHiGDy0A7aJt8O96fkHkZGHB4xM3i0t2xM1LzY3J+yu700gM1bEqoZ4UKcbpxkqU1DNpTyBpjN/
nqrqIYYRBp9Q7LfZQAGMNH7s9hITtk/BEHc+WGWIEHMOB0N3gDcWV2lZfdmXmIM8fvYZdLZ1jdo0
wQucc2dbolbUszS7TPE/hY+YG6VUjkV4EvzW9bhifOYH1cEGchMnaH7IkY/AcPrzT8+cp4vZWxNH
5Wh5jErEOYPkN2V3EfkK2h/7LhzFWaCk1jZ425MUuwMjt1tiISSFchHi58NjRAUl/Vv9htevuLCW
W9BDT1PJkbUegONrde4FdysftaySa50V/Tp1YbHK0KrCuegMCbxCKy7d+WBFfrR5k5ZOYLjTCpMB
ZnEWBU1N1HlACHBaNku/4qjVXUmBK7l/UpLDmmUC40q0YRMycHQzkicugH72u4A9NBwja+TVrwNF
JRc7/wxEiLQWgqG+xMHuN5li+RGFHJaISl68rLjUnlABrgMXJTqSZ0kyeWzEeNhQsB/5LxOLUriN
D3VTIqP9h/HVlZtCLq9NUQfyn6YMGOK2rKSq03mf/RxQSHgxVOACG4HvsjodGxJezwoxD1SASyoM
5WZ0kCixsJ05DuylYrZSdKabychcSU4gsOZOJ9Q3eYrHyEZujS8nxcz7cuhM99YyNJInWPfyzazS
fGyEt5Mhn/cy0SOeepfF4Mts0dS2Z7BL4jzXq6jcOfMXPRglEuq43MzM47T0iUrff/83xVd5XlIw
Pl082d99zDPV5YBDPt5q+pYiD0flOAgd0j7Rbl4QUrc9go2Gv+vQ5H3fMM/LN2ge2uQXn1PMAQh8
3Y2+L9XadMZ9v+kDA8rHTWXbPrzsnoxoMR7PHIaM1ZvSGXPUteq4tkiyTq/OBtehRU7yaWX9PRnN
Eb1KV2LFYW5fxBZwTP6wkFY/aduPUgC7hMBQ8Bkw0Wc3wp1qaTKodlydn9nUwZ+zMMge2e9DXwa4
Y1Y2gcTmgv0OtNBMCRPNU65eH4h5L2cVjRORb1H+CkVKPRcmqrh9wclGgTbTspXzI/fks+hNk9MY
yb0AuEGuSPOBC/5vuDT8ffdoQr9D8giqMbTVjCTl9VgZKhIRjbMG8YB9ReUVuv6poM26X56zMI4K
e0OvwVvAhAhJpgczHdBB4AwMFNKg5GkED9ipf3jaJ/Zix6lzh1ZtwuXLeNVnzDkIU/Q+KQKuAGau
qwXqeTD1XU+9RXp4UsgopH8erM0b+Uhk9Bwbv83BJEobn6+WrwmReMJDSPdL0wh9HNCWkLjR5VVx
paXxK2T3f5GVXtf7ePDgFajMQrXFQxq2mmUSRlFE1w6kc/yR2R/wsDLKWHw5RjBmJSICZr3iRgO4
7oBOLLHhsOHdJCFTdBNEMnKqCXxE7K1ERL77WnaVTkfSE6MegExnHfdiKakgsYMDo3R2Kb5wgVGf
dT0xNe3SQYBcYy7P7UdcifZ2cYJWkk84mJb1L4ukKEuwvQgT5XYY+YOZnCV0t+PY/UC7M9bgp1AX
MXFFznSmtFmFZfhWrQ7okIZYflEGxR7ZGLFJPEGpPN7dDKzAmqE7ZyXsDNQ2TcIJ0HKp3G40C3o0
yEZxopVNFV7Ko7z9dsT81B+aL/7zPt05ahdF4B+zxYZ+eZxM+BBdhEOfA7d9lkwFOvyId1GNWouK
MMrsFEsgLLAcQC4r5TjBv7SR7YRF5yDi+0BhkDKMiZImY6lavFI9+WfRemVOdEgfFshXTRBxW4HT
oY+uiixjuA69+8FYA5rAKts06Gw6O2cAwGlq5HcoTeW+H8Z+ZnQHG9vNnJWZCp8lD2pRVD+gO3m2
V4OxSPRW+Bfk2AOtFqiKV/kpLVlfU/3VqwmH3PbI4m1cEoJQCgmY//g/oJnlsG1n4dWUEfCDvWTc
U1NarUaBg2Jy+eFzhxqNvdg94L10YnzsQk6iQ+zcc+0MsThJ3OZ0cnkBl4kieZKxmQHtmeqkQbxi
yQQg0oeAlgOQ0hMC1lRr149zRjgdgxDSZ1EP/aDM3akjpWF5qSPyDFtWtKrgsgiLdv3Ir2/06NW4
gA0KXvzxt4xSLH8nLTkO9uNX2Fk24CnuFQj4nXjOYVWA9sK5XxAqHTnfeIyr3VMkmEJkgB07oNLM
h80/9zcRcDyQeWmNwlZPhMEnbI/1BkDLYj7ucTnL+5Jjopc61nU7MqPAu7k/AifOHJclWfcgrZY3
4jUbiRqXE2b5kLlyHX0+htkNVXnrji5r5Qf9PYcKb2JexSKA1UNqi1VVG/Bcj+ECvd4ZEyHiijwV
6x+UltlRsJEHwtO5Zfsou2lS70jIo+Bv1iv9MeYF9V2l4m5FJv4gTdsmDn+TafvSqTk3YF/qpJpd
Kbtb593g/kfhEwUFG2Kmv0DO7vSQVKGtJ9geu1X9sF4ysiU3K28PfC36WJoXvnnsx8mZMcDC96mT
l4LUEZiQ54BAFgYSQN1jifpUEAVur9joxyCYuVvZpRulxJgS3eS3NYHyR2l+xJpmsfEf9cCrR070
fH6SQFALC+OdJcrs9K+faNBhBQe9bF44OFoEWu7AqwAF0Pmhryb+Yzxd3FpYBXLGYq6BZA7NlAYf
WF5cPgQ6HWFTlxBO2gwNsEnbUBg7YK7mMKujLpuZpsaiFQXlLuE4kERimipRZziZ0Wfo5aCofeFT
HWYAi5nKQsvGPxtG7pr8mWOtbyb0GsIBQ5M+S7neHpXUeZZFG9pwR/gFgnPWg/K1PmOzzDG1aSP9
Qs1D6Kxc9zGobvA3nYS8et8PSH5C9Cs3Q6KqYkyVhM7ITlT0E90X3b8y7qYIp4UYP66zGkwjKWC1
FUoEKlWyWCHF3JVIsstCDgNrxcWKbJT3p2+QWgk4oNidmXqIhX7/bb50bniDiHZW38hd4MwMIHYF
WoxOOQPkgo6wweI+B6+mmnfIwPFupmpitYHBj+fu/K+VLwI7hBux9NQQ2Mqm16yZNogyeVhKwTy2
n2UqPCdmHw7B2QmN+lr6V4TjbKxROPNc3+wC7acdqcamDPoC0L0VOUE+ADb5shIRRb6Z7vdLnwsC
gUUsRJ49Td54D33Q57SZBbZVk5CzUQmNRFdlCtFua10Nr/7fBszzfKKFRGlYNjkJ3P6A1n6uPA2c
XF1zrT2I20OD4Rm38ZfB7nsZ4z/gJHKYPiN+4fRPbCUNPVWai5D3pF+KmjT3G2wDWV1iBBF9zgjl
GPC96ZysH0yU3C6zfTRUYOHmpmFrk9GDKEcuA0eKtU88d8t2XIMRAal6jjGhEjfE4yI3ym7qNqwW
4nBMK5w9WdWoAsMle4I2RhMGK+vTK/rtIjh0jpwF5krqWEPMTK5f9Aa8WVVzyW12mCn25ESomfAH
r7VWUbPrrfTk1+a04M+bW6Jx3Gd/m6f+FgkLhOrlpZm5nbeDTdQFAZCluB8upI5h7+MclF3DibE2
a58oXHNV1XPwlXEkLfs+Qwecp6KLY8ZfQu6Ck2JVu49sftj/9kJv+a9Wx3bYoX4BKFtD3FQhrWd8
gambPqbhNTnBkUYFhzE40uPBuz9g7OyS17yTHp8tIpwS1N53LfLfjC4AO5PzVD4XYfDsOI6sCoIk
DUYPQEhBNCoyv0flJUMS3GRsTOowZEnG489HcSrDVubBot+ROM/zoj4MfkWWDRKoRFNDGWz59QN+
iee33nfjzkooS/8v/MFOVvKlwo6YHC7LlRqXLYUFt+zHiCMaTl2snRVQQvQ3gcf5TKg50U1UCjD8
EA5Zajlld2st4Khy6RPV2t6lBgg2qCHJ5ZErBwLG0PMO6vRSkzY/Ug7lxUxGin/uFCZBP+YK9Nrw
m1lD9vHWezlhFJEWp/ITXBAOy5iK0hWCg09obnuvQe89fBXcME/16YYyE7vjfQsUiDqNpnSZ3yk2
C8IE9+RzEpC4rjQvkGxiVSyNMKB4Jd4dbHkqlmdGDqbXwUbxigDyJBrPJrUTD/yCbuUiSayGcfTU
IRJqRfRgCFQ/Yxm8tgnQU+sR1o0+SH73E7bNwm3e90DOxopjWzUklqIXKHnwR6LWdtAa3J/FIR7j
wfPwLxFgwCxeasVxwAQj/3lGMb4fcT18cfriSmuytaYdSeuB/+UmMb5S6foDSF6IzSxhoWyua69/
rwG4x38hkQYsPmsTjN2fIDwhuUcNzaz+h+WhVPl1hw0c+8qwZAtzx30YyM1c0jrltIt713z9uP9e
KBm/Onk0NqltpPLG4pb9zB0rJA3qKJW7GOMiitjxOoc2My9PY2g/cj3N93ZKdTJofu4eyRMEWXwa
c46va8OwAeC9OHqwdQQJ0e/ntrbvaBs7ST7xCMUDVzEg7N0sHkt1Ap32v41bcHiA2QmTz2V1mY6n
DvIkb/M3taMdaCBgBmQzTBcqjE7Zrt+K11o6u5XH4uB/AGdY3G+SChoCqwFkGYpaC1VjwpXGuu44
vufJMyNscuCya22qbSsVsPDHkx8ByAcVacwRx7g/HgaRNRIquC+nydKiLmrwLXuPGZaxLbRr8CKP
jxabew3d+9SeTanLh0mTShVODzT7oO1ioWQfkLOmKmsMqpCxyCpILXN/XrHJKlYpKpfqCsgOXaOs
Ub0lcRUym+3b5U+nY/ZoLOvpjNRUPfxWBru4ZBSzE9b7uTuRIIH0dMg7jLAeZEQmbnRshUxigbVi
b0OUrIZBLeF3E/4ohHt/UvqMoODIxPQWObBFWBkqil7oacn0C1kg6bAuJcx73LIGjPl4sKXKg4Jg
p3P2chHaZZFbWLWtXKGr+92vH/kHI9UbgBx/2g4x56jFhtpjb4GYdB/OZ+vIlgpRcBrH7oBaSz79
azQe0zWnAJI5/yOuU4uRhybDs6q7HMrc2t3S6vZA4tj87wXjbhELNbg+3GfRTNQ8pD4n78wd23E+
2/qKy/elLgHV/iK5o3QDKGDWesK6fsxtjBYDlRgSsx0fFPaBjkQXg94TptkT2gCxqu6tfFSNRQab
EIhN1gahxA7J4wBoxt/uUJ2DlhXtZVyOhufykudG/7FUroqMkvKFsYgi7TEXeQLJTIT37N6XAR8x
H7WCPncj/UjQFGsCVVXpbD87SBwXBWxvJHjYtpL5KWtzdo64rdTLrPc8DBEKVkq5iuuJETxYGr61
vy+dfGy/aIVP88uZ19B9xh8Ug1chKIbdUk+gfD7QGWpkusW7XvIKht2n5Hr2MhFxfoV8mJB+B8XC
TfJgDqIwC0iwKUzCo1nYIZnl6yKjwbCN7w8YUCb+XBsmENK3wxJuGU9oawCIdvRhqtsxfR+qhKIt
EHppQ03ad1hcmzuq7WYxcx/O4J0l/BbjA+3x592ULi2DThE6tlYTHm2N5fj3yUI7Efyzcy15Mh0x
xJOfnpmeLFbpuOz4EI3YNpZGeEicSll346neJZouN/v6yLiAxmcIDTluC4PsW4R8Rv7IR4kah65O
kQgeTUCP6Venh4o0auZeKJvp8+/AzkY22+oA0HPbxZimhWPibKShJ2VOLcbzwuow1Wb751cBCAne
lMS/v7IQq1VcM0jylaIlmPKtjTiB3cFqrPFkaPb0ht7q+QhA5goaPnLZoyKEYxQTbLZjlk1sfHLy
MUOq87SrgDzT5eA545fWmLojtSgbUoefMuKekpsSrCgHfdn7wecfJ8DWL7DEmatQARE0GuEPB4xw
Ue61ipguQaaj3AErEFJvEqtuJCG+Vy+tMfxn/SYmB64TDMeASmOE1S3OfeSzbC42DZaVd7wJfnVa
oL4TbRi74/satE+2g1QM9vgEJ5aLTL3f1OZsV4FEWVIm32MHkgoAxBJXik/YE29zA5diZIAaAUSl
dEhDqZ95rBLoGcGDB0Lm6jK2/q5GGvBlzNG3XFvr0MU06IG+zI/1XOghGPU4wwO2ZftN08dGUt5A
BupwwFmeWbWJ5tKBQKIF8+MvJEQceuPSpUUl7jsS1/ENoEAg61gutDmFFT9uW5JnJ5W5gaxnp8+a
5b19YzZvvmf86hsQtmdneckOHDrMVnLF6E51IULUcb7WxA52aSH/wu+uBGyDgMmjQj0Sv63jdbiu
YaXwFcBYVmgl8uogbfsa6YKJkFKdpR+cW0f5wqcDgk3yC/e2NbiC1v3WajPoY1j2Bm1zcbcsJ6J6
Bd8SExMZ6B2fTDeRHpPnlYZ1RisTXgjFUl+K465waSUELEuNeFmpKLUf9dOha88XiHLxJqk0u7L2
ZekQSrmEfOUZaW6eCrDH1DPBFoR6Z5WQEvyfGUryyAIIq5L+HVrS66hzXE8D3N5ps+/jVurCWYvs
ePB+S8oBve1Wfvpo+TVpTSsuVX5u2di3rrRvLP+UyvEBjZ7bId8HwOeWaxZS6x5IJxi8fU7UsUGm
yiwCWn5ZY8gFPmxfEhiOlAgPkgXW+z/S8KaQ1f6kpwzZFaTzAVsUiucdOshfnhkG276DpWoeugJ0
fyqGGMSOvuckKlWxBo4L2sJRRHpIW7039SvJmLVKC+5QcAo75QceHADiB4CFdh4mTL6X3zTshYCk
gfwljvJn3uGVyu0xiLIkHqZBLK3nokqkqiEKb/zXYDMHSsoeyAU/Fg+femQnNZGWC7N2CFwKGlL5
hiKxOOXit5cjikf4A5hFbuSG5wIBSZogylniX732mojN4hPuUb4vPArkgeqNDjDvTs6jPu6v1+L9
8CjjA+Z5Q/E4Hx9pi+dc9pkM0a07az0xocotgrR3fr/2pymGnlqFVIgDjDjlhCYaBzp9v3qbx/Cc
5cu4SBThIO/JkzPW7kFWwRg+oTMiamWQJyzSHsGljufl5CtpN4aNYrGM9NXiHCirxf/2p56zBvGV
MpRcraCW3mEu8klTc0h3pDikYJImNTivAUcVpVdX/jw2OKSBap/g26ekAHa4pReKlFc7AFSbFJQ5
Hm/lOO62rG4nIAD6qhLIHV2C/XufV/QxEDbOIUModp6bUnM7Tw+S8C/NTW05Ff3ipqWBqKoQMNGD
GGmVU63qsl/rkKDXmmzWVyFo1LX3we1zyFYcvEiaFDgdH1kMZWh4f991EfEjeFbWxad1CW8IkzXR
m2bHzhZpTx+LEuQ4BW1pomQ1lcutKzapQcsdScydX0WOEID/6U5SNvGelN1ppRg8wPMcE+LJZ9A5
eQws+zolQViVOzVCs88lVxB7h8eRhHwhkqJWhJXDTQI7xcpCmYMqXCp7ZfJjvXx/1JDRQJklPQSm
KGxgi//KxgqyCgF53aHqg3vH4zuFIgffUGo5Kal9kD8oWBzVrWd+AzpQCalKxSWzpN5h06W0VtOB
xC3h7p665qwMVP6TAA8uBKWzcveNYCbOqz9nBiNJdlDI9o7l8ZFGRhLc2rw8dKs4e6nnShh/KUcy
Q46zv3aai2A0J2g36HBm8jymtR6yH5PFP4xRmZ5IdFj23WK+1DO1J78tiyOi6e1EQRjruyhQeT5o
m4CMzdsTOP2eixSfgV5vz+xr3VraLOKs0edNO44l92qNaJUgDoZqwEsFNxa555op5bADR6UVoWYE
CC4DHfOtWBV7xUexHPbbIu3++mO+7W0ptKjrXJPpGPlgBADQ2d/wJ6mTMqr0lYBs7Kb0r1ks/Af5
WPK4hp+xZB+hB30mHxaTwvKNnYs8ldvxw1Wc0k+6rve5z0dzulwPyaPPWLGDEG4vwMG3UdNsw4KJ
UuAtQpDXUAHhlS42WAgSWbF+LVlDjZ7ohfFZGeGj2gxJTmAS1zAgFPVj9w/jPSlb7rZ3HuBlzdeM
tSnfSPtbcsuYPR79682XAsO9IsOPxL203J/lIRlm9N6RAK6BZnV5NnWgtVpAAaDjy1zyKmkkDq9m
sQpr543wKGvMJU0Q8YdkKwMLWFhcV68GCLEeQUjWsPwNyfvsZFhvEJ2lrRjW/18TBbz5C+JgY9Ml
AqVMmqg+//pOn/Tog51sjmdWT+gbtSnDbDQyKX/YrbFeThVi585zxtlCso8sW8+bu03oDXoLHsyh
vUDPEkRC4bcPAHrHOo63QbPUuMfZNIZV0SBFklZ/P/9jbiMQ4bBHzv9Dx2p155JbfiqWgV9Wae1x
BSe2urAPfPV4ZzJTYDYEwpkKtoFpK7cf1IB21JKZl4dTZpO0A46v6Xor9zSb1GNcCtzD5cSTIfN+
CWoMUuvCe9jqnK7RtVKkN6Sh2f7gGMYo5jfnLjrw33PZ2GJfoXAkbh/wqn5NbmG2HHt4ZjKbD+N9
PNx6LQDVx6jOBhw8BEc/rjq6t+mcbvMrVLO7rFHlvyloaL52H5At4v1eQ5pXltU/dO4zp1rYHjni
6dVCE43iZIyo3Y6dP0W+W426R+NFk9R+Q703Xrjsy6KwjpDXYnK0MtXpf11zJRRIz4g5M8ahCvK6
bmv3Epnd169nuIf4OSEpBNOj82FJuwcFYFwl5BLyErrw75lo6FYR38I1JNNMa6vC8QDoGdtM3Ot8
F9QoLdW0WbR+D092QxwahERHzQ+RPOEsAPKroaDiYsDgRnOBsvswH9G8FBc86o1LjAtaAcVtGbkZ
9ba2GnjDGOY95cslRaU8t/Y8p+r0P03tF53+VODfj5zAM7M6QVhVFVH4EN09dfotPFZ1Rp+R0ttr
7UbdGBgBoUue9Zav4KRb1xc8JVKVySB6q/nYX5KUcz4/uqAFevcVnBvbg6qFJckqnQoIip8BsQ2U
zWncScCosQ7VxzYWNn+5s2s4SA2vD/RiYkk6D+fHedVaI/c97nkrnFNpm/eirtABJVE6pcBNg6uM
GGbVK0/IxwQKT3eudgRxybSTz219gibD9HAbpzRCZcZNndT6dI4bvoZzfn9YmzdWvtcdrvmXozjS
u3Ikhys4GrpFLMGTRHzVjedKMwCnszo6yVfn7sKW9S4ioe/YlQHyVrD3Cey/nEoPplFezxEqfBqV
aNALD6RR+21ySGFwmLs5pQfB+1af8WrLaiwH12PFDiv8RItit4qsNMUNxhAi2wXU/PYdOb3STaZL
223Vege7YrhDTolRtnSJylsxgrkd3cbQTCWntBlf4pcr/7WGTHMrokHGIQRteO+b3X7GmFTqSJAI
+xe0jHhDDsYUaBu6xOVlB0s2vjbbku9K1SOsx6zTw0vxZIu7cwloHEyS0xK+KPlFXN+tcc3beqrS
Qu+NmSK/UQBwiQQwZu3BzFhLDhf0nHl+ABksv/V0jLlIhNC0n4pnTqLmLL+SrmU9uEP+7TIeD+aJ
pkuoCRcjAOVIbUbSTKkMgbuFBzMsaOg2TGT2byi1Ffa2vTgalICzcN0faKqeopd+kqwpfmxjXJMR
nJ8N5S8tvBJAOJ+BbJwTfbbsEFgJk3S71HoZGZ+2ju23RM8g7DholuRFc786mW+CbRw/qypecHxC
JEgp8gkMv16UK6BJI6IaCzyZUyBruF5x5i9IlUW4A9EsXAI/mBlbHgbSVaiyvavtWY8TE7lEIE4L
vwV2Zg1zCDATpZVifjQJRY5NHqqGRS1GfaOPpegFEFrer0s6k1br1wjpoOONgANjkkxeljZLP8fK
kiL4KWzj0ao7nblSO+YtkrbfYouRj6EV8Ga1D56QjlBSvSamEhYTDaHy6e5MD5bhCzB+adSI1RLE
CkfkNGuZjjdSspXYUEhNFDdUMsZjwss3AQktCHqPiSulRrXv/qJQuacWC5X/6YiDW253fNNQ9G6L
11CG0sg8T992YqdnH0BzATX9JCCPcxcM8HXAO18gNUAoB34NB9rFO0QaJVq75KX2rBKp6zIGBXvT
aTZqHVJsemo25exy/pdOammI6Ry4pF6pfTN7D2UYZVWKpRDgWvG71tMrIMXbegnDaJ03tNqw5U/a
3SS+UYXfYMwpR//OYYXzARXNDey5ntY1YTKzsO//7ryyRfLVAS6kptdm/sQ2eYApXh8NrWFbuc+c
/hR+YsW0cbU/XpCkD8Lju2VWWriR6IXloqQ/VOn5f6Q+9XVsKF3seXh4tGxsI90ty3h3sir3QtmL
mlQ68z0AgF3sayT9fl3Aty8LSNEs2g2vHBrEqAID4R20nP/o6P22RI96rv0XMnDNBxM+nXtLnQWT
TqdEzqzmvNIC6/wzt48od/cgv4mv/ZEz0bO6O8Ic8DASfic31odC5gp0e1jYdTNmFQ5V82nX1kaW
xL82KIjb6JMHBHuBBbVK/GIO+My1vVbKSWQsbF7CGd/xEa3ZBBXIpbgKpgjI+QnW8CQd0rIf+mum
kJ9eotv9AHDHSAMjDAOtmJL/0FjtKVbUZQlzKRqAv3Sb/cRWC4vn11b98wVgRanLIj5J8CtbiAYz
ODmhKpIFANKMLh0HDDai5GmaVxkf8Td820yf8T6PJgSH2+Eg2QSRhVpLyDBBDkSXaRDWoEX/7dOa
3GUzmGMi8W+qPrXxaFGQaguRyOj1M4jf53cJpKirDglrZqzaAAUwAmqACT41yD5QEo6qB/f2l1gN
rEuwIgmTGuWJJ54PGqtGCOXgHC4kSlIuJIVfD8GJ2nGmAJMK09CEsMWYwhlb8ZYqsf1VUsAr84uX
WtMpemOgZjTZYZYU5e5iWaauNghxP6eDFGITzPagEp2K53q37ZCqpDDwVCoFLMvcVcTNPoLSIMae
jXJY3QDVr/9DDuvCk1FhQsKkufGePUj7ednhrPh6ggv7oD4Jy1hH4ZO3Wpe5fwbcGaTRONzQwaFJ
LIP33KFeuFtvYmr6HA4PuC6qfvgwApOWecUjcnIBlNTuAI5geTsm3BmFjIaIsjsd9ROPGvJh8Lsn
vR31VhSNyy3AmrP2bH4/rE06IAFJjU7t04n5hMzJCf5bW291ArbEeJNL9xoLmIOsr0T1R9PW76PG
4l635gf38OC3+ggkJsPVJE+3yEMOCPudw9F7jU767+P1SrkqZlawsXz1rcHauIl9f3WQdY5TJNuN
th+ZcNAMyAAj7BhM3XwOuOpMquvN9Lc9kHTsivH4VUrKBRc3Q5NZ9Xkq5P8pguW+1yTcb4Dg3rdY
LJd2ZcLc2BYYR7adIzcUSY5L6BMe9R4QFFSu8wWRaaP2j7sJpQ5svN5Kdgi/hO/neRJORIizvqFc
1pzTD3hcncglOsFhBNGGuErvgSw/XPAdKD7OWH8M6ClvcxHFvFyu0eGvA5RMpPAIVMsk3k5AduWq
qElTNTa+yyAPVyTUMRNUMD4GgBUqHcM2obQnadMuHHr+MxVTVwikvEkwjv6t3tAbN0X41Ln03XZr
ufMQBLMaSeHbVULi7txlEMMpaNnB0OD9zbANTaS1RTVCsJss7tst0JOKyWXdfB1EcZFpBGMmIsQn
UqvEAiFeZG4REfEsUkKvDKFnQqUBoHY9/o1L1Xgy/3neIvIRAKFR4vAN2GpQ4W0pt4rCsDo6/M7H
M309anR//KRAQFNyCwiOpI5MmVYkN1cDTWGgOhhglsBao5fuIDVYryFxjCiUMU1CqFYu9YUTq8a+
O1RNjppIBcOpCp+zUSnu23Rwx2/kDrV9tNbCRBjnYD9UJVXoJCdR8b88gVmHWhhAlYIetHACvvtS
yHd2PSVAtvycBorWHg33GLlIxCHy8w1/X02wMauCfyifZIBsXHOZr+BtC8poqYdnliq6c8wVYtFC
ouiibJHki87TQjHHoT7e4q3GgC36EBSRhZcIbEg5CV1DYSCni4EvWL3gW/XNB5TS3glcO1LS/Mpl
RFZHtXqNbFgUv8usCYIbpTOTa1mYyR6xTxTACF5yVe8CykfixYsUrldXvYfWPyXRce/nVBdintY4
9rRzXuZO6hSCD7K2ZHIvDIsiM/rL5KKUsXe7nu7lYf/Glg/fT58nTWaSywRV4tUcVObVWcBSeM3K
3DJ687zF7VjdkAUiJYn35ze/p9TV8nB2RBwxKhtQt36qTJZHzGeN34CjcNemaTxnR7Fq+kY/yM3a
toCafqX9opWg7FvwlQxMsOoZmL/6drD8ZWtpb0e5acoZEYVeNQOSeXicvBKixGBS2dbUijOe3zqh
isODStTbEmyQ3WgqLV7p+ZDUX1ZhzeYXj2OgXXIHf8sBpyLyKGfD15rhIq0/cMfCLKKC/dF1uJXx
tBsypVwc2ahxgUJ9e8MnH9AmLwglPLOTsJCoL0/rBKjXCetP8oZdUvqkxLtMPV1Tcsay+5Fc6FWB
sEP/gFxBFuSj3mK7T0VG1PiY5o6s2EJ2mNijoSi9HT4m6R64U6eJUdu5eesGFg7Uuj0QZbQqswZs
Jh+MhDphxhnDfBItfOXZKk6qDZSoh05q4xNnhP1ZjuNDlW6bHi6gANTpQ1k+rn3X0NjW/UMK7DhA
75riB6dCfPWPaXfbl/onSf9+naoxy5zaw34NA8DVPb2U4M8Y37yk83jMS+mwqJQhgES/69DvtBS1
b6sQfm32BiumtY3bRtUr9/b4c0sd++HSk6fPsbYxA3NgAfuwkqxR1dTr94q2t/tRItSU65MN5UQw
EYm36VxB0XlGP2nro9FDrqjXgAjjYlZ7v3bORJI13RfBMzpkevtpVye2UThyurDx28SsPQJt0m4T
xPM09iR5kmxeQG2gSJhQtA4UtFB8TDa3pulU5x1b+HJCfBzT1EbE4kFZEL036FGWpl+03EnDIlEY
El88yPb6NYsKGkQjhAYzqNfPZp1BBpnH/Z2Y2FAgxbepgIXIUxSIwFNNp+bWj5pBWOen6NljmXZK
tIkxo9A0LA+ve/e7lUXOGUKmRbLWy4W9eQjExv2j1H7KZS2DLmxHgLFSn6omeHQOoi4JjX+0o1r4
xWi7o9QTKuvxu2Iya+mrXHzfcsxzLJlgeXXuADoyvmSt1ZAA6yI4cxGF2KCx+TgmVhWocCfoKCmg
5s0w9xhBG98y1TLScyBUdMJpzj7b+frEyKEgckVG8HZlcIQYnulvi2PPPKZtvtN0LfKKDYL4Zx1E
1kaoOl8Nv7maEGrQz9JKrTNjnq/EXq0lw+fNVtA5TtFgE5fIdVgHweP7DkX+ij30AI4TqLmt9VKR
k6Q98egrWTExW5WH1fcyHbwhBVhsZ7SIVOmlp+xOmF4alq0OtHXyNKbPydJ6sKpddRIwsVVVZqSD
YIVH25uJOJe6CVcLXhKwBw19L+TIeDXrsk0qJ6YRGDDzpsMxdj9KS0xbi45bPYpz7Vl+U8bwdi77
G2f3J9f0eCLIQuEOlbgxp/3Licr1Sc9K04Q0CRpqEdOoSPPpdoTLX/e36ecA52u/US2ykL71J2qf
qurmklNrcwN8YTm85h3Z7kQgwufJopH4tuTaYvzPcmzgtq52WPCi5kNPn/mWcqqsm62Fw31nIv4o
m75DLAM2u3GtdxqPc5+LvEMXwBmmnEsXpvDrNKhK2HlQTxMBpbI7IHZnSOvKxazHr37LsAfbDvbq
JUxoUIN0rHtMe0Ws+SSL7PXeiMqb0DOrupwfipkFv2LQxLNPiDJWs/JrO852aopeBgXLrWNes1Uz
QVehvMeGNCGgTl79OlUNoC7Z5mLDDZu4LKEQ9w66BEDO/ISzT5VFSGZTjn/RCx3lDdnG6fxDxxpG
XGpWBDGxMK/aEKAj9kzfo8Cji6ecwXplWw5lqQpJjLdqM/UOo3yCeo7/ogCIwTTVLHPyOBl8ZZ1j
Il2hH80oNU3eSpXL/2f1+YSXIsLxjCltESxFrqv/c+zX/0r3Dgdl7rn+ObG+am/dzAGX33Utavps
xyvu33r/9hGI9lWTjZGdW8UDyAc7zWwiOXvyNPGTlq/qqNo02GwaqxMf3KuBklbUj8qttn3wrU7u
u3MROOQ95iIXrz9dnTwLLfyxvPKcqdOVw9tn8n20vA5WCrZZJwl/8m7o7rBEl15GEzET/TeFVyQx
2EYDzRSxyOZ1WgM3DzexKWMWdtubHshR5P9zElkZDh5G2ri7JAjSTpjzt73U7zAAIqCMkLawJLRu
USmJWkg2WkjQSOLUHRk6HQ5wOrXHqgnRHKJcxMG0HJR/w8sZZZTPqENpsbV+h//L2WczzVv0o70R
UL5Y2hYlOb/Ip0wYmdmbxH69KfFEL8UHednIVg6eUXNMHKLZ0QvpZxNbxai03Z8v33UdnnMK2r68
ysEXWk8S2b3VBVoEEHLaihJ70go8hJMGXn54CXHMeaT8Wp9qcXyK7UgnR9e6pE9hOayw09rVKILb
30KOg2xpxmixpd+X+EheL4ivBlGob09Rx7shWQl0HTIzC0bsaveTBFipRjiCr66/pQru8gdbqgTN
Qxy18lZniPqdalH2M0hLW13gxQtzboYBkmWhtM6mpC3aiqNnss67eLUxjRL4JCC0uLqSo3EMffaz
cToCK0cFf/s2QTz8VCb+uJhFVHOuuz8OVDVJnhNKlL1Gq7CL1jJ5Fr7+GYtah3UrVl3lOJinViJB
qPisHORV1j0+Ljw/vTcLDr0d5tVKO4ec79W+W8kNZFMCHX8wnF0lZVOWlPsoytP3GIFiBeYnbF+g
VGybo+/RBgEQOT3yMATMMh8KMIBivT04FHBP94lK9KL3Lp0i58IjjSob7XmMf6zJjmXn8rtqDomA
Spz+r+0vJf5PrZHkkVcXMrUNWR013NDZYebSPtjMH4yctQdQnaEWV/xm7MInFDqmkI0CtHvI3gNB
bsK2wwiTis+fKknccgh/XL+aeVJjPFxBKiuOZegRvYwv3mchYhWB3SbiX+EEoFvLPU/RvT0n5SEC
RjBVHi56IeewX19XcTeK5kOJPXhc7D8UIC6LkdLWIoqrieHTeT7I8VV5vFkJYGdGc/G/OUn6Iask
Ff2KYydJlHduF9HXGxsK87Oizgpye8/QhKtThXuJbMTZBuvkDqZwYM1g5GOdr7jcJB/jJNnTnGQh
Oljq2PMGGIRwRD0YwNaVuCujLRC4yOtHMJj1ESdNailbNk871ZLnLseK783WnauaSrqyByl9RXkl
8e42MhWXrmYqhelpTxH1KN4OQNPfstS/GZszDyQ9+L2wOjurtG3aAw85XV5y4bgLgwU0xx7iy+Qn
zsSYYMkF5MzY9RsKpPjzZa0YqVubS2okXZWONl/WJaSvM8kUNZUzkDUd9bgGJ+UTYLKjRoJtFfuq
h8S/P7YZIZy1H0/nXdLiuiA3yxVJLw3RQz3KVIN4JHDggd8i+9vDLSMUEfHhDnOXyGvL3cmCXXEQ
chUDAXa6Gq5y1R22Sjx004fsiC1a70naP4j/6VVmmKZQ2tn220DZIRuJUHG4njtF5SGvPaPqw+8u
yVOwaGNmPE9SCCEKmOs0jz8RMNP54SvmgJ9f8p21pv85l2hjMGhHdEFwaULXDsE+hjZlFPERfZF3
gbZkJBc59BurYJumfZ5/7SoZcA33Qy6ur3PRYob+QYKSye+l0qwE+GWf3kjiJyTUyb/gqG1fPk4E
Gb/oIYo6r9MyTX5k2dSUOfmd1wCEkwIOHyKVVcuzkyQzs5JWhpTfuAlXu++GDUjQOTH+ko7xUj7k
1cdfPKHwm5JoSBnezcQ5syudUquLT1grGfdxQm/Q/60IIXIn8OPRohgMWsgBs9eGHZDbI9uBRKch
m3+XhdYPTSRXwudaLAX3u2nOvYqWSM/a6rw2r3COa8YNXv48yGlway0DipE/FFpO38XvnMEMenRo
36IhaDXJYMifn78JcBA3bFvXkRyMWUKttxgy1nEdt83yQnC4zAJoom3FL7qszFPvkN7lnrGtLN5S
vjU9qSwbz3TdcANCnuY4H9ojqt/6r2n6aG0a9uc8qYbQ4R/DqZXG6MWwzBLGB045bK59fH1ByAnt
8LlK9RAiH+nrp2DvGTdAxRscwhmA50qHFW0wufzAze05+pNUlH1k5c2rYBCKTHiERPTErt7Jlivc
3WhnUX8F+Ax+p/t/GtV8jd3ehfG1GFtwDMB2yTG/+DdEdDWf+yIVybCxxAbAvW+U1OY4iI+9rmAR
gAdY0miu9xrXnvGRH4MdHACatvp7nlmwz6KtW/fNyCU4XYy0xMPmIHQdmvoTutWI8s/fhfQ5CLpR
KOk9UL8Rs7A2jd48P5Wic+5phvRl85ogpw8aNeOtmUtcVErq0ekieP20erZRN+PPNRx++qxiAC8+
zRqJ3NefB4Miv3a2O3jUwdWIRClNoG2teZnyjqxZfWXUBBlebDRiF7rBoYx7lLjsEWQFVMoX2DsR
3FC5Rw7uDA4xZTgGp5yKMUS8NDhXEjEEP6JYJe3c/iitZBB9Yc/DjudFiGESgqoRCLzwSupgXxLa
emNYFpicWbjkDOacRypR7k8kcIxBGuFkGPx/zPQ0tre0kgN0JJDLqpTyyThB5OPISjBDn0hot9cn
whTPvS5jddN33HVs7/zc1f9C4QINhE4e+m/nfpfYRCXhYMLjUbvXxdEtNA1MCIz2N+XnBTxDXjCV
XQQJPYl7kiBmc9XuvxQ84wCY//pEC5WZRCcNXn9unWrzD1zX2hz6OpViC73DLGX07Z2WzD2UEfNr
jvxZ45/5Elgl9yr5Aox5sOS17UeDNZO90qdhmv1gPC8sEDjEvhMI4dh3HjCnl4fszBmxRL/CPNCV
8YnTwZi28b5niOduaYu3jazCaX32v9Ny5ZNuPUmU1olB9PBDRxyKvbBkfD6uqFcSkIiflEqjFgBG
sFJeKojZkqr2BZb4gpKbHHXxUJKWlw8wVtD2c6AhXuA9Dntb32ldrwTHUnQiHmQL5rnQKvb6QDPZ
fbZQxRmMrFjzRIwoJ1C0PnhXLx/nJXsGpdJCD+M1epcU1YIbOIeTrYvjkeLLknaNsZNZq+9lD+0J
Pi2OE6KykIFpKdqbAuHkjdm/CyhhNETLJaJM20GqzvmsnQq6MLA+ARU4IVRAYFt2v+5xX7RdIgCs
jZnx6B7nvTfT1exIf8hSn1UfzJHvLK3r45rCXq3ok43zpZQkyrQnO35QkE5JeuXC+/5olvuMXyaO
AbK9AiUmGQZQmAP18Rd/p/40xn9779C8BdRukQK0guHPZotD5vLqUsZlIlJaCPt5snrHIaz+AiZA
yLa8RJrIZg/DqWQbwm+v3par/CJBVPOOTCo1oayaEJXedRx6O18sGtQUArdt5W0mJBxKxeLTuNZg
NNVVCaggvdKik7CiggC5vzlsd0+kxXxVlsLEyWNkgpBx/rO5BIlMTHuRG3R7YwvF/O3GSCLS9uQP
b2NY2jnNIN6uZyIgh+eTWA6Lfd6aUN5FjELCCTHQlyl5wH5dDvaP+hGP/yjnC2383vmP5P6c4pOg
5O/G8gUajhQXvoghBe3wUEtAl2deM/Y2tHGhYYOjov1DBUPUOHjR0ESFXaF/bkr8ivC3LBR42/hL
ZfUb2dRrrFNHeMhxaNG1VUkY4vIsD9jNIodRTmQQdmibOUzeF267YGGjbPvvuyrY6J90YPnKkBDj
z1YcLbPCy3n/WcvqaysYNhzods6wbvutriJ0p3IstKUTjSMViw06BICmvD02BsgM2/J/uOJubc4T
NqtYA1p53jvyuJCNqm2VRDLiDTUP5/xxn544NkCN2xAELJ+Y16XlUM9T+CRiICimPrLGdo5XCznJ
EHRZ4TLdwxOpjnH7Dmas2n/oew9EbRe30jyNjo+pkgME3i2xs/sXSM5TJG/BIMipkG1Fb9DppQLa
7S2Zrb6x82Uc+PWM/wowfdMpBZN+g3uQB6n8pJsEIEJfGpW243rOmX3z0xpeOpfHHi0YxAFflsET
4I8aMLl8jeemHNX8pW+WbkY8hBjJsfq7Abc5G7S5LQ69soBH/DYtjuodvsGrkC9WRdU0U8aXkcar
QSp5Gx0lcSK5pWAbD+93pXklEcLXcqh137Ua3JkNP7ELxgP9k5k0vZZWJCy2WhWaPGR9//ACGlNB
AHElGTOeoSASVt98lEbgu4zYyAbINURxIzktgndOcBVjJUZERkBNZxIb4gB5GdRoP+b3LhFliyX3
Qw0n8tZFbfNbbG81+xM5UVEFO570QOVC07GUw0QPX7pKBEP0B2N9InkD/MXV0DTh4NK88omw3B6Y
yTFVmfPGvxgmxY/tDfzsWTT0DBOPs4RaDQDbHDmPr9QPF8RN00067RgAPjaS6ApJ/nqXbMcOTppr
9s2GLgyfgMHUwYjt1rynREjsYUiGJ86Al02Jsld9zhESvE6Sbf+qaBqvQ6/5GQPWtj+DAX/JveMv
eHOZl1T6udgVfj9f0burEoW9j9KRethulaHwkESyPkuPdJ1eWH9VWEBkeTHgvJSHYCvR8fLTyZRG
zgZTtF9shd8qBq+rMYxrEA4gedNcdBno9gK7tupS7WhWUF/kU9bGCdUnAG7b/ON+CuFDdttRSIVa
PXVc9g4FEEj46bL6J8I4QXH3RxeWLCknfe7iQCMeT/kIQYUtNiu/MO3YnehGQWUZ68e5N+kj56tC
HWa1kDhWtD7wYL5vD3uPGzBE4guSZSBes43LEJSZyW4wjFW8ws/HuZHCvv2oVVbGmdUnph8yogk8
B9azdxVP2DyYXqD06sClRzBnlIxUabRrdZ9lML19xWyWGh5yT8tGmJ6wUzFy1NTi/36GOp61HnSR
+N0jrXAHz5LS3eWEqnq0SXUmjJ7YNYvGGL78WqOUA54GV4kZIlht4pGRhNK6Nb3+b4SNf9hlCPv3
Q1i1imayEs8XMxaGltkAFnCo/CkaqBOVL7rTh8mtrmSicAMrglhP3E5L93Nq+n2ip/ZNWYS02Og9
Q+B/KaOgay4twsE2VSte3teqfWISbFJlt9+0UiRGlfL8v/PYlSYeILoa+BlHvC+YsZvEr0eIBuqb
UfObOvx8tOg+9046Q9FvZVl1oDbf/8bJGm91Pzn2hjt8CDac+18aSarSjcAIjNm97jnSH0qzpXcK
ve9hmWI9lbdR7hW32nArf0jFLt8c+27XC0hSTkZnWWMKuSsx7/NQjH7vg9rI0DhFZooPLTosVwnY
j+Vt+XvrDESeTlSpuuqyP4JlRKmQb0YIuDR+5r2OQbmqaw8I13i9Wh5Yr5CdH2AfS+Grazspl+Yy
vKD7UHrSLtTDVV9j+faHvFJiplzi8cPb6BuLhwkQdJ5RFH6L1Rvtb+FHsE7ewHp0JIlicJDBrdfo
jiMTGX8ZFRfj0XwDZFZvykaNgSAYD/IRb/H997bNt+cCdebeM5+YTZ2dZs8zta5cYu6l1NnyZvZJ
D887GfUW2zMgU5dsK6urRd1VM1DfUR6tXX4RHw9uzwo8M1fVX0QXXVi1y3GUK2PxDjmWX3xJ9Hhx
2fXK2HZkZlXlfrhRtCCsHUpwyvL2oZ+haaPoSiL7iSjWazk8az2tkY+KbBFwtPU/vbIIA4OKK+P5
GbIhqLF/gZg5z7zdgSStSGOwknljaVpCd+KGZII1ilk6Ezr4DK3wDOk+QaWbR1WbdTpQcDN+fWl/
zVHyj90gi5TYA8Qke44j6XjDsZ25mlLiZAj65DZFykjycQKrHeZvWYuefyLMEBLhWNqOyNDzjaG4
/c1xq636J/LG+8HWhaXBX8AN1kGLuuAJZK23IZvfqeemd915ltJ8Kj/FkaAnCfWLDL4UzGyCIgYZ
5c+W7pT7ixuRQE6apn1W/qC4UpsatjhMqKy95IydZDn6KYDU2jH8ijZhtySHnnZd1GqYgHQcL5Qq
jg65sCAOU9cWbLt+7ZhdmCcp/If1KJ25UrstrTCyXYiWuyQoigX11zbluk0r9DDTVjES+GiT1cH+
Yb6F9BmmPKoxL3RKWBTi4tnCs3MIaG/4U/mTDbT17LeXr++jfWTrHMA+N/hohqFsGRR8OVcTzWdB
DHaH3O1L3tWPVoQ7GbBTbxQ3lWnuV2Vt2pCrD2pecv2iGdK4//rVOFWv/7zSVtfDk+uILFxbOvO+
wyR/ELN3ta/hnK4P3ODSn7zXdvFMCpgHXfk7r2OkpQSCTFPpmxfx85oNH+mCU7zgFk38QFFs6Gx8
dSv0gcfpAmRXnB9T5ukv1A0LBRMIWgQM4qyZ39CMML/U6SmLbA5Q89AI512iX+9YnRYfH0VBWiwB
v+HwJcQHsrZwlobIzZxxYB92MpgSv5rhjtPnln+m3fEPVPbxSWpRsE7j+5iyzjWQTjh0s5RlmXC9
ocefXIlX0kJi+27DZO1w5cVkT5TQM0EOViDumiW4qKdFE2WUt5S1DTCWOTSGsWL2+jn+EXszkn/H
aZfi0uf/eCa9pKhsNF/4jzY7Qn01kk0jGlkxqvCN53Mw7OaseBOGMV8jsJjEdfN4PzNo8CsNWOKh
0xaISrbGy8JhtY0DWk1CQKIqeWWDYSEiZXXjtYgaLLrzjGJIW4yArQFqvgvdhlAeTIYVvaOql3uZ
RbrnUc7tKCrHw8iAvSmgzQlQWcyVm0gnfbyMkrAHusvmdvTkfkkOYt+9aPYz8DXZ6Xa23cGbayCk
8lGsqGy6XqN4kcqVgbPcbIDC9Uz05TC1HFhuuzDR3guOcGhGzGJWesXIpInCMJB9nbU0M7AkU+bM
0sWHQXx2ZsvsySuZEf38LZzsIXNcMPCLYP9Ho3YnGzytZwVoRVvzNLuKtpvqZDXogyavmjZRIXAe
XXDPsV+8PGr3h1pvHMbGrArwJXcvjPatkZcV5y+OO35r1uzK34xgq208BHJhHJ3a+bKFMgHX4b3f
UZ/MJCRWTsmJC6CA7PnC+WLzwrfE0aidwvtQJlvCpN8rYvj6IcrH+wZ1oDYZB18b8zbrrq96XQBE
wmJYKeUjjQyh8kq/SKK84f9nNVanTig9VhYX+/RYDc+wbYs7aK9BLUnObmvWq/cFrXip+Axqez1i
f8eWd5yzpXvHp1yTBT8l8sYicJuKG0R0glFjAJUWYd/XUJlnSovP3+27ysipnxnNLYln1p4Q/SK1
S2/ak1DI4pNzvZrGv7gNV5A+L3kGB17zsWMyGhSTThATR7SQS4LLUd7WSbDAiKzhkE2bo4Z2pZ6P
+azdp3AQTe/ILp4H5z9kKjHKTof6ZVHADvkmIimLj8Aur2ABDeTiejSMKMtiAhyn/tOwaPhdi4Lb
0C3oJQW5GSupTEAmdptI77Jq7lSJ8SI0c1gohu19p1t/vXcFAB0iOFh/WYKL606er8ShxvLfNFiy
2dQmigNmrbXWcVtLD/4l60VHOQ/to/JSnV0KXEYNk80A1IDXl/++2nclDWoX1NYBXgCBKMWLAkMl
gWwUG+ielo3sHlL402ZYBTGLNALlYDrgNVfPEKS9rU9wLMFLXrXhmYGyUPilh7ykGWgaPN8eNNGQ
0X/rjSj81X4lNau/gJQMXJtXE7tggoG3WUFzsQmk4IaO9tZkf6V5SGKhIc4+w97kXsF5yzAIt0eD
Bw+tBPI/cg787VtWdAKlCrbZOfK3jYoUmtxGIXrzGCkl5ivBLfiC6LrO0NxKVpkK30j8ByMsWhu0
FNht5e0lwx2AmP1dmaMEKhPBLcOgAryrLW4hJkq2FiLIl9YmGIjJumUrxdctZq39FoNaOKFx8d4U
IcyLp1LorpD0oPOymilZg3OPc+53kCMIchu/cugCPywxLH7QbdyzNaBVfr72T1IPG0xmttT4dzlc
UkQme3ByIpQ5y40lwYO6BbnhYJ6OLlcoSOr2SE7KZNWgEbPzJ0z1ezEv2o8WF3vlnR1gZTo8zyN3
vXFTKINHo4GXpDB+qTTfL50/v0AX6aT1NPGkc0thEU5uMxmoMj4+bdX7JLBWYhoSjXPRcjFdw+1/
ZctySvZdOEr2BZOhv0O4k1SlW8iYfYtq241h8zwiEcCQoHOI9YezvQrbFvSH22iNWU/jDAKub9rz
dsjbMBn7bZFAiayTsWiUgeQyBxFjf+3r7G4ZlabyRhvTCpLgetkV46+DgTWu3S0foancSVOOSgdr
R4K7Tzv0SbDSao558sHsf60Vrl/JVWpsDNK5RDEJaLfW6xRt4lsdvNVyMQIYhqXPB80MaouY/WHB
jFirpvSXJ40haZV1dXkMxkbV9M1ukU8xwm5svAGpC5dLo8FRocQFOoKL6CNTnfPhizsdEKZ5j9SJ
z5bHG9EczS5FeodupxGt2puCRcIRh+UQJX5Y8yvnYdzC6mTITGYf7IAf7utJhE0mObGKeh1+fmEu
mkAbif/ZNaSDwbpQnzSgw+ebxt8pEToJjQfcIQKV/q8D2KZL04QLBeigZ6MNJuz/4CIFDpw+e00K
tTwhOWd/CjbjgErpv31ezzPsFml1HJ+ra0kaSgsX2DZPIPtPm2K+KY4TJ6HEBHHp8i+1EaFUdvR1
PRxhC7MG7zvSqWzwKXrVrSZjh0W7GfKSpekU0Ld7aWvk3TlXoRgBZDKfW3GZR4Qq8H54AgqaUIO+
wvde8C0NgWAb/d07jeJJDIlKcXIMxboKTax6txwgtaDDcGivlLkOSxY4bsq5tdQ8cMFUV3bVYg/g
tMxf1JL01bZlyD3L71lUj8Xi/tDEQMH9+X26GdpJhP9S2TGt6QPPyUPo4qJ+Crd8fzCxTvIZX2Ad
HiCjy1qKi8ZTnQ6lY0OplTdI10pNkwiqukF9axgMKy0CKvQ3v5MI21Crvm0QBw/inYmtmyr3nm7x
s44EJ6Jr/0455JW08x5GXvFjylvgPUyZ3zDNULPGFicK2y84kRxT3rXPjCgEnvSWLT0/bXliMcoM
yoX5LTsjvOhKlVQIOlYrnyKmnourdBBMMpM2LeDF0PNiKouZdq5LlAwnz94B9FURbi7MoeHnONYo
BPDdgN+LqQ4jvCaUcDtG/NDcd/MvWVR734izGHAbkoyHlaih65QOCJmNsNV+ZUyOg1ozf140qQ7P
laPU70HfpsKEh928R6p9h+1XzZCHc+zZix10pgbUCxoz2D1l3EVcLZOhJkX/JDEkoe3xYnBXxkE3
yhpEO1gDTnBkqzqC6XgQk16OhTBjFsP/pwXAJWm7xwKPfNdePo+8FEeR/+3uV/v4MkxXsD2FxCDk
ax4FVQXCuP1CksNEGma+UNscqd+4fmuKNfuVBfe7rol4lc7UUDxemi52Ap8Jer98sYWqYthDjYVa
aBNyZaPpibuPtAvA1TjxI/wII3QfQsr2PGnZATsDM+uk5QB4KlrSlN/Q19eaAqckuuI236VcWB4r
LsJmvWeaetDN7AUJh93p8qaBunvlwKMmad9MreDnsxE1gwEDkyOWe5Ef5kdVoNkZeRfem6Y9AmQF
ne3a4uB9jOIsAEKQx74plO3RfsgcABblzikJC4bJ/3naPYQ5LvQzuWccIVYtUI+xFBUXDId9SH49
kPj93zFtFWe6T+EoXj3gxkmcayOAnC/UJMfWY2VF73j+uNQ1527hb8jJt6pVj7ioc8Ctmg1jtoay
5CD6KBpV2zvnymcu5Asgyv6j5Ntl2kJ9R33PXjR0yYw5c1ZC4FSXIfGNwKwkueZLVqchGmGWNJyA
sS5vyM/Ng83TawHaWVfbyvp7M7ll5zUsGZnl3QAk4D5qSrhMqo3wHa9rM08V5Pt0EQoXs+jQgQJf
UVnqLgDk9Td8aacZQLkH0UQgqY4h0GsMyjAi+YipszBJGUGTvcl/bMyWtfgbN6fVfSmn0mlgOD08
pQ/7WV04CN79cFOazCDAJC3UpL22HZcXh97g52AdR+RShBPxTnm4uacdYhBflIs/y5UDJvZWPeka
0zMnKiBu7VHfUTBT4YHQE7ZlB/L4L+WlkEwAHfzEGS08cPzj1IAqrHIil5kfHbJ4EB3qMVIcMy/T
ako4kleIm2p0wTolHaG3h0t1JsISTAWVVgrdDV3hyMUAB0de9YwbMtDl6ef15qRaWoyz2rJi/+Av
LZJeB1Gq1aj75LkoMzPEp53RPHhm6xWfhu1XeO96LqehClyiaTKcULU7HsG729DOnb7NtW9qyZ5I
KBHr+P9Nyefh4aOB6aKFX0jKDL5RLqHmqKQg1bnLX0UMr3VDtRfeglUSBgu9C1+nbixClBGHj4+u
qpB7MCOYqG58MIW6buY6vjkCg5CoJeq0SoDuP/8d1JIF21ZWd6LsznBq0Wn48bMERfindQRPbRM5
59eTV49dt8iyYIkD9O4IPk3fFfUd25OkOL8r4og9wKd5gSqUD3/wshsDZyuC9Ci9Cg8XkmLk/85S
gNFhJga2UZWQlpym7IVfqVl06OIRiieJG0FeocPBbBKotnya4wCZAD8J7oI5Q8SQjRnvC74t05QR
nsoLxp8kebos1wNiIR/zPhG3yDMQnCtW2v4eKuBpT8GgWvQWFu3XJmjGNthrl8roJ4z2tnuv+tsD
DSpmdVuzxlBxeEIB7EjPeXreeWLPgCk39ALU0UXtOCtqxsSaGafOGxsPvINLIo7lFrpe72rn9+in
v4ujvql7prnh50S2c8jf2pn9SWqK3YYCFPPrT74+7Lono0eWqYxAbc54VzTJXzkDn1YdGkC2JQO+
wsiEJUECXA5DP4ZZ8ivrGouMlrCryA7/gsvd72lwCxjLluVJNfVnzpkXTCnrnVX0Ejqq/Xr60blE
M1O3VPgUQdMUiBlHp6cVgBBVFO4KooZSzwsfCkAA5OXi65oZABCeJel0a8AjhEHFXrNgy/FwYiOb
jBM6ND+51uJKlTMQTAFrfDeNr9wEeloT1qiai1ZKdvk8R7gzYmppsvgapEKxyuNl9OFQEaMWtPua
bFW4z6Ku4xfAHo7nOKJU5GwO3nt+AN7hc4sBXKHeXTOlqNHDzUx+XpH3O6GhW1zpvgC7+cEueFhd
wreWpleNmzLtLS+7JKQ/3kkb691UbhDjjAJYI9Bd16N7ztO5vOyq/OdJI0MTgXltKHl04I/eRxEM
rkHHg6mr94q8d45zEiWFtYrOpAJ/y9gthEKRVQkBs3XoynAAa9o/4teTG6YBUv5ONCXxtCetRf1i
KxeYbkRuXcV5jXoYPcGI2hDt/gK8kOYlHyX8NshgJEc3QhSWkiMaRwHo3wjKqQ5G/xTIoHgyc2sl
GzhTZtY9tWzQL6OZ4gY048FpwCSRF0p1Xz89NHYqGw9CFGzwNs8F+gAqYPcW+ZQBpbZfeYp1nI9S
HARTZ6gzbfMrC9wm7lbrbTsysAH0onOEAzEyz+xA9oaKbXBU86Ya5Vmfm8l0gOYT0K4smepHWhD+
ivojtHbGJdCns8eKGL2208gp6wUQXEczCxAzOmX/KNKqyGLADt23QukoqbV1aplSklzzlKQFMgVe
pPMqAszAfZuHfr0UCq6i21z7CPy9toPGRbR/QR1EEzg5cyE4it+Z3qBlyY9RmVuwU5TAuJrQXz6y
ED5XXJD52lywIoTUqk6X8KqMWpovuQ3ULDPdVsLNWUzP/Ud5zcMENlbbNBHsxOVo6qqnsNDTOTZa
KWvE1Ch/PgZfSctCNBYYHAZVQAONnxz8ALCYcHID4l4/f0N+1UHhbcCBFWreSw95E7A+mnNDGFig
T7L/RFOseajnxL+JPdhHidUKAfLxDdxikeYa2JYg14t+Jxvn4pDr+W3MpHPuoDV9X0zh7QpedGvs
EFq5eQYuF/5aYk6qqSqmjDddgyNeInsd93YH2xA5MAijaIRpTEC9Us2PCAmcUGcRClqgpRZUQB/l
pB+29AwHB0b/90g3XsftFv+W9EXaKscP1v/vik7ZNWKWTyNoItNSpgaZJTHRiUJaJgXMo+0Afi/D
Kww0Stuix7ojd5Lh2FCT7rU3LhLNZ7rwSy87gegkP/oDJa27KJw16B4b30Gjq7hV16rdTCHmvuqw
6O+EZVvi/LEY8vSx4RhGNAuUwwDgZikrBJ320T4RF8zHcpYiC0PvU3tbUQvVmzJJllQtBbhL5c6B
FaFt+QvwulrEtgCxOBIgtC7OLQy6tR87EZRMbLgEOKJWYLBmvN+ZJPyHnW1boFy5gj6a8eMsYXrF
YwU/Db8hmHDNQeGN844+pimahbfRlPs8SDmbHb7D24dzmB8Vx1DEOeIxXAyhO5ca5GL5NyoT64dD
7X5Gv6jKcN6w8GnKUoRdXiSgGleclFuhFUcrJ+LkvqFgvU3DzCw646QpW2JXArk+85TSRzbL1Cak
f2gG/NYwo9WjvgHmEiAc/+Qztaaz0O3n9/edSHp1vlZmNikfODxaqlBlx0YfVjNSobthw+T/gAQN
ziit8kzGEfFu8vvJv+ZDtcusHWQwavTjz/qWvAoPrE1FllN8ug1DDqRNumeLk5aJwcjcK/w56Lik
gWxwN8vqZaVyJKsOGvmT8TuMWC99EUeCsBuri7JbAGSRP5EMeSYVu49aNTJoo07X+W8bUi2QSm+p
7fDSwMVXU/6fpCtSjXooe20FOMq/pNoRMRUSkDv90EzHcQFqcpN0jOMhlagdx4e9Bi2buTZX13AV
4VDB3tU3i3lWFrZH3G8BX0mIbQ5H+mcTMQXc0SmRmOJB5liQfEDAqq9ETbAkDwvONxiwCum6f64I
I6GHI/wFKHqWHVyC3HA+R49rA3S714XdZU8akDs7tqsyHOG6Pdqwet0y9lWuMzaoSBD01oZJXnQd
YJXSUILunl7h5RQHLIEoYWuvwfwuDRYdyNi3h/7MPb/MKzxluFM5W8REdqSM8CTzYcFtC2J7tgIv
oUuIs+yDtdthY8b30HehBxevvxUs06Hd9fM4fWyPubUTdmGffKFaF34Kjn7x/mn1yLXY7jXzU0sv
vdIoiYuebShdQrQdRQTzKCJ1V0sy4LOfuG/kZ+V0QV1gqd+pTWh3DKbYZDS4co5OHoRnzNN7Jo/F
3VvEHgpzSbK3MSE4GuIY6KCipl7QYMugEhRrSFYIVddSXG1PbT78nLZ2DF/x7aS8I/h0cGriGyrB
DfO9KY8QljBFt8LIVCUWf/aEH7IZJlicigEA25EoFVNTfDIRzveQjIWuLHl8XDZhD8K4xQHd8EZ1
E5FjtzGllr2K9HFariWY4oN8zObGwId6/WBfCill48mISxZVnJmQ+U1aCasNiSECDI8SfIRB9VBf
qbw/B0G6QBGqC12ynkGN39HShhuOBF3ZQPQb8q2mjXPJd6jkOk2yILspDBodSsGh2lKnXIiY70Ka
kTNV615TwDzhZRLjzfFHcWyYis37wxtR73EqFAaA73cCr06l7gF0Q6mzASFHwHRbwKfGtYfGz3Rf
Q0VoGt1xfslybdKOUtHNnZA45DPTGghem2Udg0Q7r80Ia8LPGwZRvWqI+nkx4+Ix0GlMsF9I5LgJ
+XjWIDNJFWO4BgwV7t5JjtG4lBUVI5TA9ujavCtNzRzyw3Z2tG2C3aq5nxwHqwS6Ze+HbDH/p1n/
bUbmdGj8BT9463xrO0z7AH8Itc8QrfAF4vTmOWkh82Kr41oyd2daclXgxs+8Ch9h5mJfKTsJEhzY
wFi7RWE2XBMwKDcULCiOrgsa8e2eVdnhx80nVoQWvuqdGUjuj45XeceSHSMyU6TqxR/UybCj6Zqw
M93SRkKpdDHbLZGARccO91kQ9X918oT4WWN0eQP2K2i12mRF+iSa4aMZejPYVeTHNjxu8k0V4NYj
M4RGs6wl6tk2NRmPY1P3RvYI6B7UDHVa/le9vVkpIRX0tBFTC7S1RD/x0wgdkfpE0t/LuvWFbb/V
P1pSOwKXrOQjSz8XsvR4eo3D5+WHcSfy1c4PHQVwTPhk+IE5GjMD0645Mp79e802dXkEAT4Y4IFd
RsD3xp6ynpMKKoHSmsxBJuv09zzId7rVHpfteDgyHQTwv/B7dE5AKLJatpt9BHz9FrAVrZgggksP
tCCz8cj8RLjZB9M4KSVS8BBuK1vXaNvGnRL0qcT+2ZwzDXs8mYYzGVpU2hggRvRNPLblbEALJ2Kl
kQEDcJTHl/dQTLBdgNmwz+e6140LjbseWq3gASBiwUvOWzif1USKHvbozfxLqnyShmbUTJB0W4I4
QJeR1ZhFrHZk8E7hhlNjEzDeBnTZbBF3T6NgXkamvRw16xELZ/Yy726YzroOD0644HN4sSkbiwUf
wW6/zEDHLagOZq7tRS/BQskO/zbACo7zfIQ5ocFKuIynI0mld9xFHqgrqIP0KikdHcINF302WEAD
4/uzUHuYWtjm8O9GffbdBINVKCqFd1obyelnlqXc/+Xot6I2eecR8snV+F/ptrNr5UC/Iq1BqFn6
bD/IANkTKvVFh3Tfr90gtzBGa6Vm1O4sx/ciD69AAuUaJzQKqJmSql9n8rB3NGYp0VVx5ls/1zW6
cm4vycNqH740GEjOWOT3VsFTYP/m498mgrBeWKVqAHaRf7LRpNcKCiua+3gXXGo04A2hX/9koDlL
EkDtSylZ5dNJvPgSK6e2vKP26oRsYaAz8DcncYfVVymgxJK2sI0xWDEVjdSQjJP3Fz278eh586XR
h4XqB/t6BGmXEMgzBeaZh2nuI+gW8YpBqIr0pEXLESen+1bOcmY1IbCpNKeuEOqQ9bdZdLVk4RuA
2lWWe2g+rWKZEBT/+KELYXZLq9DogrtNEBTwypGjIqGafR7STtruLLP1RNWc1Ut04zsfaYo2pEPC
YALjM4S3X8r66Kn805RCTdCTJZnz/HmjbLaiNGgEebFEu301JPP3e7SMgwSWzDC9lXSSCyaqQ7Om
VTFNhpjmclTtF7so9lUDQ/vj9uk9RlaocImfnG+3OtH1x90HxDBgmCvjhJleYw+NwvmOBb/95qM2
H69VLlx42Dw6y76d7mT/nUUfePSZFx9pvF1hgR37PC+O3fA9N6YlA05sxx7jXDaxNxrxxC4JZl4D
yQNMX3DlZeyv9BVYpL0H5OVtlJFIRROzUghuFEUqUzGge6alnhrid6q4s3xU+7KKVtXG5UoKmR0Z
R/lngDW9DyYudXpDcsZg6jYPMZ2r0V4obPQupyLHCRh4B7vZijDoK0WKCZ2FmCTqrcuhSXfNK4/E
V4b4RRbEsST583L1Pt4/OuxD1pfqBk4SByjuvWt+cNnUsAH1clQK1rMIQVE2z5LMkdWuB6OUywIc
k6XyjSaWXhWfrDFvw42WkyQESu5xEnn9CV8vKJ2RvMrFckfLojVfeQAicCX8LPlsh9IsR0MRGfvP
jM5fL/ZtKXD0D1HLMxiMqsV/Zs6vnlMZ+6msL6QRdYw7iXJhQQ6qhGoF8W7aYTlSkpROrXQje5Xd
6T4wOyVRsu5cL/If7XsxsDafl4WhFTqBA+h71k0JiHvk15FjPPUvS9m11Tq0Q5jxj8noGMc2Vlir
zbjIgdHbkrBcshU4D1NIpuS4F56J8Q7Xbrqe3gMI3SLbnolXqh63DPl56MpmHAxB0q6LGn4AVLeI
fFIBvn9kDZ3FeDFpWB+EQvJJ14/VKBcOLS2Mt+IUaxJAy1Yu+3Nwnh9IgnXaf4RqrkL2kHHa3ji2
RVoxTtlsstnfNB+e19spWRH+WK5TUU02wOuQoGjofxQPjAdMQGkmoaGsrAACh/wt40wo/H08c32n
oj5WSCNP9EKL1STSze/adF40GJ5KVDPtaZM8pJiEEUYjAVHm6ZEJdi2j7i1HQpiqpyRN9aCw5XJR
1a1m8I1Hp8TnQkt/UzsQYmnXruIq3rPiV0CQHR/UcOyR3vyyGggnrugD/fAJtj3j5evmqcLfqlou
+6OrFeeTyd0K+x9RMSt11BzOwaULBi5827oG0j0XbhEdmgr2FjZ5bGW3CLeIDT8mzw+zf95q1Jef
j7tkKk+NB7Btmq1+d262Ru1qwCYLAfluMrpVKROVYHnMMLnXOY/AEwnL1iuQxxKDb+1DH1a1PpGu
wbY7g21gTmI5tY2fd/sZrxBmiJz5Sj+b9GhpUoFcqphOncfyYHYscg87jAxHlPfdWvdkCRQoa2Ze
kdv1F+mD2S/tBbXdbGkzpK0KUat5yhOK4KTYcDNRg8CBKDqWQeGLk6gX39iSJpdPKd/CfHLxI4N+
lMcSfhcrs9ssDdBzko1ICRQa3yks8fwQ0HaN3xk0o901klZ7e1Cgpc3a2xwRowlUuJYdSstX47ch
+78Oh6RuTSoRZDEhz61Em45nMLX3fS8ZL509Onv4wyPwWFMwVMCyHi+csZThr9zdaQMNW8vWoysQ
lnBT7Y81HeHDFzN4jT3YYzGHcjIkkmUGQIJxCybMbX220BiGEFr8RG3s9MK3CKB/wzePX7Mb+qWL
ASZCWLJm+zpQmdvlvrYaM1FMP7vEHzfGalzeKlIG15v/sFlY8WUYBHOT7Ku7H4DA+RPHgwC4tv8p
xwEfK5lTN+3ImF3w2aM48jtrfyt9QJb35Fu1ApYcM94IlgThBer1bpLImfCQMk7jciVzq0T7HtNh
eXYcFMP2PXKmPKyFLYzgwafBLvvfSvXdGnhI2yies6KsQwQWkargtsu5DJlVeL7U1k8jhAz0KFmO
gtu4zVn1/tkS0EdinALRKsKD4FOcbHnCuPvExLHaiNAWbZ/a2SImLj0UJaGBiZJX5/SChw8WbQoL
78nKYRwYdQb3rtDd79kcZTkgncWGZf6s1VOVWvnfaokWgjKI6bCVi76en4Ohnq61yD72d6xOeUku
6HkMev0k0qtu2TGisi7UkZDHiG5zZENGrzWNMQwVbTRdbbA811tSAUR7kjjrRSLFThM7SzHKJDgR
1tq3vr9VA94XnCmoIEiCqaIunGNracIl3bzD6OpNhav2o4gpyg6PFgkbSRqJHRdHB+egM3OLgoOT
BVnq46qGMSwzZzqeOsrUchWSAUFLeddFLoGlyjaZEy36jJxESrhMVzJ2CXN0x5ExR7xszmXUgiVu
wSzwXsNKMQdCPD798SLZu2Qn2NSURKV2c5InZOf1bPLo76elyNzov+yvOpe7cYKqEPkWE9XMDSWH
ZenqfwQHgJ1Wrrcor1ezbsGh0LA3x1Ek3FiKDo3nLby93WDKokcXtsuqkBGDMmaBriCNpfpjKgM/
2UO/ejZdBn9xEJju3r2sPJKeRl8KvvMh1foARKYv6sKs8x4kCestmErTKzGxWnh3ZIIcbrKL53yt
y5RoioqaNaRcA6JsPMwuHkA/T+fif+kGfQFmt10b5yfHEgJb4UrklgwGZcvKg1k5TRdPnejardo3
kiUMJinLmxGqFU/yTiH6c+Da6Ns2moRUmHgrH0jcQO7WWSdiR/M0mQ4tWHaMN71GUkGtjiTX+6EM
ZzuKoQez52yugHZ0eNi54w21vQWSzi339T6wdN8p+AXvExXFlxooTTKOf6EF6d9BDZUrk+4X++y9
YooH4eS8L/wtb3uc4JFGs96Ep247UYJl7SHv1TToet413NQIiEV4oLDyaWWBjQWbwcEdVoR0bEBl
xEbUUjSov90D1qHiooIrHpBBTxGdurcdEF54d5fVUUDkAuSsEpxtGlQbfrSXm6u4vPsT414Lpez0
Vt/qGyvAEEp769YLwbWVX29pHLntmD4s8CriigVfA2LquoRN8Jcb09mdPUKn+Z8wfVLaZMzFeOjW
dK6rwwmKFKLcesq6aiPbXuws2+HbCWnQfYe787e8qnjpHKV2qfaRQkXul7LIaWdkTMB7cAbL/3qW
C2CmMNG1WBiOw9pOzpz6sAlzAjz51TBn3p3uOUfuA4hY2MmD/SxKmIjidpqYbqUsVq1PcF9fZ8up
uoQQfIEqpotDwpmfw72tX7JiHWQC4BgeGsuCUIvRA282qPysjSYkrSp+Pi6JAwEA7Iud4Zm+0sMl
DiuFIe28LVRt0Y3KdTj4820EN6CzSJEg/MVvn04TxadxEVlWv9jpjUvHhmxY6tXUJwIFsBJJJivt
QEGkO7eGdeVZ46FtOs0X0NmK1glgLdLTU/jjb7U05NpCckReOrdnJ+1On3pox/dMq4w9D3l4YQHS
eBuGBEM3J7W4zKfU2vBgjc6SfYxWss0oLam7xwjzglS8PFvo7nTFF0PkNk/iqFssgcugdkt9qdqk
A/rXVDAoyP9LINtUIkYxrzM6MCVHCzef8Pcr3bz15saJA+nP6Y1bUEU7s0FO+PEmeL/qimK8tj2G
oRmFaklloS8CipliAx7XkkfJskFWG3hUDVJYqienVN4hTwN2IZdSVteY93TwvTN58JZKT5GlK7WC
yTUWgLWoEzwVMEeQemsunh+dh7nFo6GF24Hx9NKnTZ6Z79GXQ0qNhayxEJF4phFs19wctAeVpRHh
QtnO+nU9P5aN1zMAPq1PeFGHKpuJjR6OyakzX8tlVZA66x1aY45P3109845jzzUtwTprAI1fMkjo
NMNcWq8C3C9YN6IeWQSkMuUgnoA6JAsOPAIpv/ngm9ICwc31y0rJENM0qkYwWbzzhcRC2GjSsKMg
dqH508+ztw8Q1D3Hd+ta7qsNoQ+TuIPnoOGUs6ybEhCLku+gAz/+LgGUFllaVTabl2TRahhjfLhl
RwfJ/VUZOJjFghYnmA1XRtgHITif/NCEPae5x/N+xwtJH+meRltod995EtmcTFD1nXmgc29uXjom
agNY4lqwuKuRHQBv5mzpht7kUOsC7iqQmiFtcszkcZFs7yCtLtUfbwKrH4DtlzmRXOadeLpfXmqb
0D2b7kqU02sXjhmBS0yh1CgoewjNh19TNs4reiBFWtOke18T/3EFCIDTMZ/Eo1/kbct6vuVdELco
1fZNb8JBnUZzkWrSliaDZtUqrU4yxvqIg/a9DU957552WE0Nma43WBb+i+M2PsSICLW2nIHye94D
PbiPPxYJYWvfFQ1XA4ftBvFv67zfjFO6mh92BpuWOa7smVxsVQdRE8xKWdjiFJYPEFRTiDImirGm
PdpS8WLjBjOad2mrZs0uwpLQOllMdQFtGizAAEjqHLvJ9UapQB9ANWHdqW0YbP2+NQdRR2HyTKXb
T/8R6FF5tGDd4Kuu7q1bVZkzMPYPmEjh1bZgjnWEjFXE6cchf9on5TNyJJPmJLjX/wslCT4uLBF7
OT1x4XDL2zZdUqsues420LwA/IMq/2CBO1RD0icC/6erE5DKCgs3y9zV4uxPycjz5+QFa+IgVJCt
Cug+KmqS70xCwjZEMqeop0hxkFeCCr7b1m76GwWVrw0F2mpKcMkbKaUDgBlQu4AJLT4OKdK8ZRw+
dkcyoKZ8LDO+LUpKXojD+lwrKoM+3CrZj6aaPhGhP2GMMsiQsi+iyLKeGJnBRb803vCp3dVE8XUQ
/8qUAVA=
`protect end_protected
