`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NRZcYSus3Hqh8Lt7O1HvnshMqsPUIDvTP5IO5R73Eyba5Kbk48nV85m7hlvmGYxGO0k0CjVRjGsT
W713YSpsIg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LXwwVo3ugwZbnxTTpe7twgUjxq5pPMg2vjNoxF0eyc4M6Fp0bbnAhbIRcYO/WgUWlRqWs2yeMjaj
/Xi70e6s1pK21Rq+59B4J95Z5H1ORikPCh6ufkgkD8UCiHIoxyy12rUPJXRun/mK6GupsHfEzrZh
IanyaJ2F82U9h2nSheE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fXxg6w6ZL+RqtJjmC/HllNvio4aQJ8rUPsuSW9WBrpwVzMoUt00H4+eSeiBEiQHqbki74j7yHi05
hUVj34JVwbUS9tAKYBuB/NmRubChTQ7eijN7tw8Q1OFM+rqGFUeCweSQUNRVYfffFHqCzSsvRhx0
SDEXwBfdSvjBj1ReYuYtcLpnQ/uxt14DOvcB7CSBpo8TXpCRV7FVvJoKQladZReHLrCfqJRAvmeF
/ptViCrUY5itsfEZg7Ja0SuQu9UpnXtnpHG1b30VcGjihPmXJwAIZUvAN4BsOiPW4YzFU0WovHpg
VAyv/k3XgnQMgr4SmoN9dLCPdPhWz8R9nOqvWw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iRjvlN4jcbN7WNgC9vZzODmkHbhz792IlB7iKkW+XaW/irtOLhtY6XWqqZQkL6g0K1ww/dWf+3yd
/qllasdWugEzH0rfyFo2FF266sY5+c361J3F00tO777yZwyUUiuEa32D4gpddizsJ7yLfDzInZ1t
lxpL7wNN+xcwFS6LoHVTHavlB95P2Abrn1Ns1uNZ+5HgOMnkJCV6RyV6afTHNSXHvByWkMZeXNuH
ysklx1qZv8wi7ibbkMVYN6qrWfmvvCucS+gLWi0U+8bR7l3YFVBNFIFxZNfQIU+rjTKubyMgF1+R
3MU6Zyr4jhb7SnPPWyw9IlURCcqEfGRFaFDuuw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ob3GkK5/tYzcx1TsuAIwRIdXKSG193BmKwyIepyqEYdTFZghmrtZHKrtyVNgk6GkdiZYpevhdoMA
SGxPlzABcYOp3pSe7fC9Wk/RjnVqQG0RIdBCLli/gfDpzFSeaZMCUaVStApNlRgrzMmh5wHDVo8c
9DvbY5tPYqB+brrErCgWOjW3/dqpfNvenroGNqXG0zF5+epKfGBEmeOugKxh84yKkRITBfu3bfQ8
lOD5Yc5ixmhqH1x0CuxSALBsmpuq/loOW4i9IGt+6c9BY4SlwKhQ5pLubbVmY9mCAATx+WKHfxmk
OvtDGcw9y7uIfiWZqVV9obmevO42abGjVP2cWw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b3vK60gaJKulrIDIqNGqNBm3xMWveqK0FnsmsuKkCbuc4VyR9eA5Pcg8xfqBBWC1bcct1S93Ls+o
rixNIWp3fN7uqRCN/NyrudX7fNeztrdgwoL9PFvYGuVonYJeyc71ClF0hpsirptXuhFE1uwm4r8P
wMuMf2uj3YyzxsdD/gw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
d7Lw1dBiJt/KzwB3Rw0Uoj1XWC7VrRwy2I7xT4OnNvKJ+FadUv4SnQf2od/xfmFrOAzT5au9KqUI
R+iu9moHXno1R8m91aiSA4crYAlZgQ2Er3m2vRgd0rejUjezekcLGckWg50Drl6KQC5GFcPZk7nw
QgQ/wlWAmnxVO0BM06WEbRC4pKL3/OZHaiT0ZLEP4QRUImBcVCE4gKGUMZeV3F7U2G8UGaKmjyl/
TEeDdEYjHC95S3jQoZZPSQFW0BChE6IqH6mjOHkk/Okc10PYvPYH83Fh+Ag6ckasAVv9sg/gN6ay
lYYXvbYoM/1TcfJFR2O87w7MS5X/IAdrlVWBZg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125824)
`protect data_block
YkQnkcowx1GRgaKQCoaX1FCl3lQebWHzaWMLZAdL2aUreT73OQVT2e7yez4jj/I+EIsBXmQvg5zA
EO9HygxW2G0O3Ls/2CfyAlkaYshAnS/a6399Q4vIqxm+iQKMlC61oawdTLaaXV+3M5kub7q6VD0g
eJh8Y4dR8cLBnBUGyWei3KosozGwRBKZ0USsHx6SoWMx77ULhqAge2JKAOJmQkNfaWGlYm2r74ag
VluzhKhWrylFwx5ihqJqLAS1yWPIiw4eKFpL3lMcXHf3xMOwWDSZQOnhOKb5i/2TKm2ZEUgH6OqY
4KtIy3kUI/s+mCM8X7g7j9obMiTG+D73imc4VR8xMAU07B7kidMVssSgNuPwgdodrLEImR+C0hY5
Co8paVVhiQ84mLot3aPvssntzfhbkuFghWXZH5zblkMq30yxxyN6fryj5VGHo5dgAFKISHvfUbTs
6vzAAfi8E8U1fx3qZv+FK5oMO2fL8+Uo+Lc4sKZWR18B6wIIMPhiYWXnG91DW3ndR4urzoGYH3Z+
lV/Hr1+U+JlbUAbvezU2jfMx6gbEdpCwUUQTh6S3hvhAT3cmu6uCxo89dMwdTVF3SZjE8REsK6Lp
YR+UyfJ4BSkUP6bnqb9v0F22R8ACVLEiCeETwqRBLF57xYSwvPXDs2E6XDoXDZH7sf5jdJZWYGx2
4h8l/MVKcgTHWOncsYddiOgtMbxWAPcRChRaxifZVvXK5tw85Qq21bMgO//vo6sl3iLvYEk5/+O7
1nMB6szmJ40rEh3wl1uEAhlZYkcVZ8CNELp/patIIHc2QYPO8NPA1fXscm34vtkeqMxsYfbWYDie
GB8gNy5JXoRqFaOQoOED5Kjp1W6sZMtnerQW/usZGU7R37NriCDs8Qi7ljZJULJBVM55O2OcphfT
d4lqvKpV5FAYvZAGWq6SCdgmTp9c2j9tABoSBDyPScrtWHtJn4v01nA0b+boaBckwgM94AxXAtol
DvQ8yO8yVP/ob2tlvnMDK/wkAbUb1dLITsjA5C2FmxaQmO1ztMkl2RgORUq3HXloEUfTkY3Ru11U
+g5XEMO36XgRdvgouNWuMEupLxpW5YXNAVfxIgcYORsSGF6agJ8zzbQzpFTrpbJSV/Z/mij8kB/+
YDtTRg+t0LQ0wElAybGE4Kg5YPu5hRdLC0JwW9/T6FhyjPbLaNC9Rv7JHLK4eGev2AT0llhBwQof
cyUtCDHQkx4xTcHFv+17xrIviBEqRJ9RAR5pSQtGnTB5bkZQZOjcxbvaEvZDrklkDJ400R6N+gzB
xhOatipyZ3m0uyFArEUE/ZUVuCJNCJR3UO04W814RsjN6A9nb/xhd6qtsPv/DXPw0hhdrQ1osFTm
dXZ2KAqMkg9MHF7kRLJ5EfJoxXr7rMX0jo6EAON4Q1Xiea1zg1lmK60W6xdzOIcQbmltQdDshNo4
uWZSGo5zQFo0HP6wj4qhqV6dQ+WhQQ0CmJsImJMPVbeDBwlwnWBd9+fEX5H0sGjeoPW160v1yOlD
M65ltMVBqmWVfGc0+gsE6kVQIjj1thu/U9dYgQUGiydtCst0mXFP0VYdfTiBW9Y1CfztT+Cox+5P
ZvIDwYZzMAAWrGXbpv3VoeT/pfssooxMh/qb0wea3fN288sBVijRwEA2C1S5gz+UtqaouykDW7+Z
YnuCL3vucafnfMD3Df0xKoBJLsFWn8R/PQzJvcDCqQIr+M0Tptsq29tNoCDCfj+oVRbwnByqB2Nj
v5bP6esLtyaUmDe1vsFaizSSz+ML4fPvdr4cmWZHnTk8uL0HFfPixwWRZKZuHwIQ9e1dC7kwTNT6
44tRLrNZ4pGsiIf8Jv6VGv+EJfb+Y8Z8SzzxeLIY5x+LRxbqohSkT4EwowXQqz5kTukHbYLuvQ81
Gq7zlgNnBB0x7ld1LIyXzEOUbgeTnFBN4W7UFXfC+P3jt4A7rxS5+XEU351dNeNodPGdOgaukslg
Lrsz3SU071xJKVqD7TrjSE9rq0IFw9sjtNs9ZOzYAVR5OIr9j4RdLIAd8WeeZIKuXNOxYTwNjWR2
urHaVHtnvZFodK/xsSpdclo5/95QS+UIIGUyNL0tXA8e9i/aQb99Z4DAm2a9BSK8o/wNRoZXjwB/
/eVxiIDwrxRrSJ9rvY8ORccLG9qKBW52KZmQIdDbcghb+WRl4AVnWNKgPAq3sbDAaQAXgB9ZXeCa
E7Fy/Y92P7gdMoDZghf6gLODbCCIG/LXuJNVX9vEvoBw/wWUA/ORC1aN7PjTZDOah3I9p/pdJeVu
obJZ44tln72YHN2rSbBAN2k6T/Ztal17pgvANhu69x2SnFocS0th5sKBMUnPZSQqoVC0ITG7KxAy
snAzAdcRx1j2TLNyX7vcKq1F3v7T3oxQO/+qpd5Qttybowl+DR7mHJPAE6jaWGgn6SFIwVyEJ2q+
2krFQR7zhiL6hKPTulgK1xtLaGXH6tR+1sH2hQzudnYAS0nR8+WIuBWOyV/y0/rvG1MaVKnGTONp
Qy3ZM9fdeJ6qwOleKBhqKaubN7zS4oK9UDeFWS34OOJfFQu0YXzyRsiWB7oAW7E3CkeCwMosG8+z
tOHqcCrDIjOmfwwFbp3USz+IImrcVOUePBXTD/wk9Cg7gP2PVMkzNlOfafqou/jKdHxo4+sofOcG
BymsQFlRGWJFmCyqDbhzkcovqnRsKeZIr/SxdSHUcPkHCrHd/Y3Ihz1NU1M7Yg07EVCUrX0DsbpB
G02RYMd8TwZBD6BDpF39X+zyfHMQu/NDpSz0yQFDVbvYVXHkk392QYjJI2OvypNbFLPk7TR32oTz
tdEsHyUIyEupbeBUEO8nVfbbdWbLv1rwPdRvzjgAnYrid3e4rqeSh/SxWIZMLUhv+h5/dVt6uO3l
jJNPFPznuAx9ZVZwI7AoODV2Xa3Vl4w1FZufiA1zK8G8egs9F1t07reChVLIjbf8JKbGYgrsbv9k
yjVNHQMQsLeSsRCCBhVUX6ceYct5RfW1EWucSxTjaubU2IiMyO1yrAtVANrrerKKsRwVBCCPjPip
0CNQ2WOS14b6+vTKdOvVri0loIX4fcAsT7QUrpremMKNso/FkjH3mK2nOL+0WbeZrPVqEHnQKcv+
rFd7E+rBu59KRTuyxTkS7C43SacJQbXZuxeoE1RvoBj0ziYmRfho508AdIVt5zEns90danSD9Q0B
yKfV/idmNGR+gWB5Ydpkxw/ImsBVuuaaei+kv/GmqCN6rTRjS7uO4HNjeQbZ1oMLs0rFoUJYSkm0
cIoEF7o4P0e0qkns2E4YQUfPCCZinGLGjRf7ewQTEFmiIGj48piwkRKLzW00HOMN3nijA0VTC4a8
g9FYac1BCUtRPuOh9DuQUuQKxVGSUQwUxo4j3HA+ToSA6CQg+ygPhdEzmMhXUSxaOw7uk3Eo7E+r
garxHvY+UDnFG+ZT162DLu8zYdJmMk0t+LQ2uATgJfiYO85TgcF1GsObRhyU6JNm36UITrDdLVCt
+jbTuDtsejlID0kkNNuJHKmoCFfVDxtPfdcKvIVTzILZ7jQIbyYhrItMZqYSjslaD6yEa7SxBUJL
j6O+l/hMtnxMI+yMTm1EvO19CbT7mAq0PjWStKIC4s1t5mZv5uBjadUI2gTKvBtH/Ik4QlauFOZa
6UbS77iXuehYl8ZyTeqi+CcAOFPE88XXOnbzPC9B6gsl/sv+HSz4Bnb6wVoOzy04tMIFq9QaLBjG
oKkEzhoZvSaBb2K9LyzQdYbUNXbc6pglh9scXPq9MqPUGU6A8qqdhA8ciwcDqD6ogig4GGTwsI+d
UaooBRbyUI/68JZmaEmCsc9tiB/JDqZ90Pbu5BP//mUkYKV7wm8s9yeJnpVqLUEyJHgJn94Zxp9v
VVYtpeY8MhfYHpgdk55yWvGCW6PLvxQ/yY2yaz9N6/r6/ay0NGgbXa5k1lFLUMLZR4CkkKcPHMIM
SB4vftzrS0ISMy5TBi8ZH6JD21EqPmJ+Wdhck+885hUi79OCq/GQF6y/140jfSxN0+MN379z6+y+
I7z1IOlXmDEK69K0dibFw8RXYR6B0A5NAlQbjuWKRKXDZ5y8nMxmfvfD1r+LTb595Q9LaBXDX1zZ
eB15HZ35U9W+oasHHhRqHu8vZen9fZYzREgXuD6HmKZVdtBabML9fe/N4X7W73agHtj6a2jPnp2/
AMv1P+YvscFM2ubRq8lwPN6Rbn3nNxPvlWyRIlmTc1V5NFv7AgLWIQ5JGKQjwpw3v7synuYGYplB
lVrdi1w/mIr/PfvekycSt0aVmYYltTZfzmAGgIhYpts25iFfCOTas5dpDgfOsKLhFeb1md/3yib3
Nqg5o5e68rDh34AtOElx80RnEJ2LB8wPouverT6UiIshdAiMCUi41rq7DXbEB/pKjEtKkdHwPsob
rI7mjfTHSNgp0XOF+m0arWzQXrxWrJ9vDrL/gT7AzIyx38ejI6Sm21EscH1d18rsXU/TSaEJ4olM
p6YUQBQIEAX/sNv62KuWiUxPbE7I4xvfNQ3ZK2yRiOavV21BcNnip8uu4BFVPvg5XDUMmL0NZqh7
ucR0FHwEhuisc6X33FwMv/RF8wKDNcykjFTvgJB9t1nG79eOW9rY/luxdktWSOYU1NhZFRTYxV72
flVRWdYVcxYZcL22TonZy+AJkSATzcoI8QUGROPSD5NpyX6fYuo+Tb+/4S2jjBjG8shA9rNu9Htv
Edh+5QLwGEjUMEYKWI8Zg0f5jRmId9zDea+V+ec7Vmstg7tKJPb3YRkTIX/6kGlrcZFkB07AdQtV
iTXle+kLejbl211OVtYO3TLj5I1/sTuVsH/oHUNPykadtChXJrlkzwivvDLAHijCFPdBG8Z0LY5O
P0gDTUk29+Qs3eGDZnqdYljCXL1wF/WfqyGl0QuP2L5TOyUnwfP0f7Ja08v5MLp5id/5hJVybhOZ
XbdSKOgo5LNU7pOq48uDDwPLoeNgBelFhIeggkRw6EYLTvMmIfqrw7pWILW/MqEbwHiz639zL+5B
Kk5gqVrC4dUywJG5SKA+GwdX8kRvRURxA82pfFkbI5Ecw+n6uvl5wEQGOnLJ4/QTa4SFWXnr0KF2
XSwxBbR8zAO8uZ9OSQVgP4F/roujJJFXhH0UyDaHyf/uab7GHvQOvpvQa+cYkBuxNupnhMve/kKa
Ugl9EMFxQTw92xLfMkRMdKStrOwjNBiNm3RPj74nICV2lVt6d6Twnup/IT/Vh473HJU8IH4fXMk8
RHDZPYGLlGQpnSVxmLEWbk0ljK/89lkPLNOe/QHPQZXgH/KcZLT+YsM3A+Gtr/dQQDdgfQJVMczD
EG4b+SLJ2VXlmAlGpQpfQaX+gzMFICrAMRTf7IbUVcC+ThFh85oqTGsOY3Cq5tEvx15cptafxuBA
a0SK3hBYUMUwnKAy5IMw0dyLgy2LVg+YB5CE4GP48+fjsgN1CXPsJOYDWqfDFF5PWGbAi8XtbycL
I96zsl4LKJwBVdVZPQSVv/4T7FxnkS5SZMGGzhyZLB1KbdDJju26wNejcCyHdj4mtFBSeTHHnWBm
tlEZewvcGHvJYIKkI8rc4HMJET0myNildknvl4dUK5r5OXyprHdHjaPMaW/07dJNW53AGg1K9qrs
147WXMK7WaKj2/Sd8bStD7R35NDzOHi5pqfZGmUp/pU28vCFBg9rcs51VvzNKIoVqBWI/CiuCubh
f7E+wXMDkuJPdpe8vB3g4xmZREx72C8E7prs4Z3ZaSwpfyhqrc4O0KDz4iHmE6PtZI9BkRY9DSOO
dXkTibsYwp3uuVs7+U+uevDR7Hy/fawGoX5hFkS+E4wa2tyykn/AWNCDRhjj5tE6Rd0fu9+Bsi4F
4g7aTjfTMvilgYRDnno3G73DpOHeYKcAYkE/9P7x/vFzy4I9R6u6eaRWhfPf+sVqjS/MATmlDBO4
K+1ghfA1Ht5nqztAfELWNqIz4lL1leSM1SYw00sy/KyhRwCqu44wf7Vb/C3Nh0oWQZqzdl/WPif0
EzSKEINvS50rWbBskBmj/28CFE4Z790Z10fuF0R8OMBqTQUnpyGNEgq4wP4b55qwzd4H0HJ2eiqx
Nu+9y7Jj22tq+23Eege05CloyN/HqYxQmdtcd6mXCm7iFmd16Y/1PJwoeO/apuQDBw4J6a7oUQc2
XXjhJYNxn/cu033ojLMiR71NDyqlAgpABOrod9H0BtIZUQraoQAfBn7O6T4RNoSGUoY+PfEutyQF
4WpIOH33K0oXjM4Hr52eUr3dSlEAzdqACCpdb5ZRAPTKYhnxFX8NQWDOlVHlqSlpUSg9udhLK4/h
TdZ9WFIWBQ4CLrRh2ULLP5trey55zP9DLBRzmZxsZv1WEPFVJXMGQaQB3ixKYm8J9GzhRXHxOsEr
Ld31AVj1HMIzGTTDS5ayNWNMe+zTgBBfGSeR4+/lLL1RKHk0UqSyY2Nq7E+eyI9Yh6hWRaNWq113
mzLGWs9Y01q9zUnuzLcsTA/4YQkUItrMEkYKDur9MygtTLr+LaQiSXcmcrFldCVZ/du2UmYplMh8
8cJpNWznNiMTrLrgTGn3XaD4UN1B1ogs27oTVu97fnWuXvnzwF2CSLt/+L2MrYWta2G+CWjL4i5a
Au6JgvWQPuNC2vCba0Hv4HIYMXCdUvE9W8z0eF0UI6QmYGu3Wu7MQRrIFDwDQR6wmjIr/+ISG9wK
meB2MxP6gbsll/etktoToehWWdNpkCLpwaaPGr8H6TW4U3XFm5rIGsbrMaGdT39XsxM5yd9kZRNO
s6jwfWtBuReHTDe3/quxs90daQGEDPjpP1sfdWt3/BHOrmf8JYEsjuZNgePkhORQOnymKpSITv+m
PslEaj4/uSdFuvgOkZ9+Lvm8gU0ssm9OpbpvoymLttWOU2LTw1WVnfvS0B4JFlEa4BSN/PAGjTNf
YJs3xVsHzLteu1MaNJjeIYNbFtJyTGR2jcNq9A8Ymi4AspnFWnRwrRRUeq49RfT6+vPT/EOpEpwc
jHUw+B+ohHG/6vGXqHdil2wJ+wHmvruCjd6/momRSTzlFjvw3kaq7H14tG2WhjjEOTunVqZqC+yM
zt5Nod9gNoWb84MAR6GFCf07TXTVl1KrAjcC3dTmedLu5EKvuUfiY2HQS2T7yiURdx/Nk/rC0nX0
GvDfQeW7h987AlakWEzODlP33EUnAJiWnw1XnuuWqTNwr3bsNto9RQpjkY3OCDGWJp0YNYea2Ied
kDqzPUaN4xybgqfpN3rOcG0e/Vit14XGhDo8H23yG5sSPVq0MKO40QqCWt3wEgo5i884riU+YteJ
JYR7QbFb0sZ9zgmaZQqg3rCQNdfP2Xf9iJeiGPow1Ppo481L34tg82NLppVtcJl0lbMDUvkQb4n8
FotX5FdvRpIs2HLTFxuMMbczREM/ChuAFEx4lXHa7hSXfaTkRxsyYe4E1C2umwM0rlzj3k2r018f
gwp+LGcerOCcBL9Be1ETXrEel4qYV42KEkRhjO444unYk27RVMjlzrTAX453sCdG4wi24qVdYiFZ
2fROwkt17GcXcsReqXsJ58+SRKz/U2VplcxuzQcSq25VXQPjkaRXvfeXE9TLj6lyZlw12HJht7wW
lhotRpemjCSLfopLMcARQsjXSelpeTB2tf5umabUIwyOngA3MXaS2jbqcuRZLO8TFFQTOSm1LVQY
oOReQW3D8/twyEER9rQH9NqH+Ojo8igCZsAg1yAs7k36+hAp1fst2K0UgRPFE2doYIx/alJWtNEJ
cdeCeBWsOAltgYIjBtHTfbb4LiLIRxCYafTGsIDjAq9jdn3c/p0hpEGloAcxyp3oUewyzibRDAdF
b1xCGjzn91PeomeATwp/aVobVMRX1zw/HXFw11S6BS/vH1NoKWKRrs1xwuuElBebd5IXwY/RNIr0
MTtQEnY5MuUepfVi7doZzVk3cOK/WwvFK+DEAfSLH0QgAn2tjE7ZYqlbgGjKLIysdeeleduYOyOp
wvfg3Q0wPv7bSjvltu67FpC/taTl4+ngzaG9al76yY2svTilyqWVxeAlsdlwauRa0TMcsWQDTUPH
JS5rzDDudqg2hOb6icTzN4floRkXyFAiIuWkeGIwtWzH48N+iHZ9gpck8Obp9xC5cL7E2bDxpg0o
ggLTeOBLQzH659nwFHwut8eLCsEt/42/KGnWAMBenTmcSFqeJvv9HDX30UV21G2VLXlha0Pm+4Vk
lh1aG3NyCwBjbWvsTVnMo6lcRRQabmjVwfi1y+A0Wgw/Sp200GbLmukrmocbQmr7rksFfcUnRsKx
1dvhkal/LHiioEU1sbE/5bp4WD4b89Pod/dEl2WAUmUiTXLnnrl2yJfLtiPlVMWN8D0blLaf0zmX
J/Wcmn7r4+jbjIOLS1GUM9J65F9UPbpYKAXH+R+I+7rNou2OKF/kl18es9sQ2rnc0XdscTJerLde
NGTpnr6aYMTxIwC0K2hcPZXzFdWSue9Y3wNB8rtyBfBRVWmL5+84zAm3Sknhqs/xXPbe4Y0aS1WR
8mVZp85XDpK+MmMjiYisBuBQa5JdHXTA1QKxn2xlfAVf62XhNg7+3DbwBmQqwKa8AJV8fuTGcZvA
Ax+Ii4ytxtye0ynbOPHxGlr6vL4oQ577we7P8vI+/ITCPLZrGLrCOHRcbiRoNzAJ2EtPwgmNmBoR
9ef9gLocbnqATmUUDoGNVSfTLN5d1K0vc104HHVRvsUeLvB00b8AiI6bp92/V1aOLayhONmhLgXw
aJoz15ruADqp6EGu149VS5zXzscKkSpbtMEkKR4fZxr9k8EQKREs8tTHcoljB4d7OTnTzWn9ZljH
oW0Nep3GoYboidFRB5ryMP8Uj4mcjFLcJpgK3eQnlw5htlBB1PzrGEBs2rabh0yagLBbTb5K1JSc
RDAIGzTkzo2sjDcgnC6xul1VyRj7/QqFStaBisgihbu5V7Sr1v6SUPbEz9nrrkGRJ+MkS8TULgnD
43qBepeU1bj93hIxy6fJz1hD1h/f5t7WIrU5JfEkZmxLcX3hfzmDHj4OHdyyOPmY9DnJ7fuDsBIH
jxSh55uJr9CDpkPnBkHCVYzeZKP/XBM3FClxEaY54oPh1j9A/EmOqojyteo8zAelKVs0zS2krkzY
DaAHVeMX8Vn3MOlSlhGyI9K78DvB1ekR4C6qoZtr7MFgd5+k72JkABy+hKIIVuh0opHbkpnp6gWE
Lo3MYSa49dJMqZ4Ng6QGjfIBu+YCJyVnvBbPkS2ji3S1wJqwJUnJZiPIgTdaKqqVFr+6NpO5hkqG
ArjMgx1yr4+c/H64nwCyD5fj3nHXxOHoNPNKGxDDKinWMq099hz56/eIkQQnr/B4zocNVjHlJhLA
IQjJ1PDf+IsV4YfGsq/vIy5Ff1fkDk9MpshOW02QAkcg3Doky+M5/ftM8lGNqrzV/oTarkVaLOW3
n3/axtaMxkkZlNkvXfoJl/3PEst+o9zHDi7W/u8eyofmqy81RKm564ajOzcNQbn/TjqhSsiE3HWs
6bAYl5XoMq8uHdXAEi5uqqqbGMekE7bsB1KYmGsfuWG3K0sXq5MK+ejMGpO5t4pNkyJoU+QBK44o
tyB4vc9lRKClC7mBqNO21ZHWJ+iMSwTHVBT0nAh9ndPXAW2fHeL69Cs1cToKpeH7Vo2OXELwD+jA
6CxyMYtlneXWTLcGdP4cCL105DWFakQQQVNYyYo91pF1OcaxVmatv21ZcNWsyOQ+wUaacfLL9/bb
sOVVqjxWTRmI8+jhNLAqVFlL2VwpARe8sOezT9WpWOiL5NTo+c3Iw2qi57orJaLt/lCKtzmPVvGJ
o+SN3mCr7g7KsgunMNUgmpqrIFCJIneeCAeoUz/YhMWNfSE2Os4R1lbYXXfltG2g6/yHG42MO+q6
onA20I2hDeSlB0ZLg9fkrReR+hgG+CuIIXsNUnFkwKQdv1nGj2DzYiSRk0Q8Jd0wlbvQbTjBSAgG
xXyoEougO+WXupaO2xr3wZr3EO813xJFvneqJTLgk9uTKknolZuCxPKQqQgNVQTohcH0GTzSrMHs
TEQGImVa0EIBffxRNvwb6lV4wD3C9o8fxRVxSpkAHgcPRuEVCOTKjvFv9ynA6Lpp90WkqX/AnsUN
PCqeef3WyO3Qox9hujsJ3aRhFNvusvAjyozmjSccoBz2gLCFied0nhCp8e6oELr5nrTPECCKfdv1
o9KMFJCGg5A6BytqeVnKteTTRXW1nbmQ6C8DL+1m8lfRArV4Pl0dtDPSfmGly3blPHUHiUIY48hX
iIlTVkQ7triyJcywQjQjcwOucgIpiqpQLvVhajkKnbw1EaZd78fwYcChPhhpPArNON9dnUGgOqKf
356rzBGM9gX1nahPtsiV61kXSPXi0DUHfFp78hg0cOlEX/rMukNrtp+HtDtoO3RfOJ+wnrnFmRFl
AFxK5akD5+hZWn7IqLiLwhCZ+cvM4+iWbZDpmWl2WVGg7zY9dLJJf5IR4uq+bfJCGi4cdlDdmZBA
tSKzFEgZo0TDG8O6EH3QjPKN/uyfDh4gnyL/YQAizNl8zPMEv5ahk7CrjAiVISSX0x6o3NPSRErV
hbtPi0UBcow3Jfigu7t9UxnrJv7RAAWyqFC+ilJCvSldQYvikaly2lXZwmUG/cIRcNvwXEanGUWE
0WZOCRGxbg1UCBx3Wi/sSsi9zSv7Vto+Udyp2hOuRs5GcdT+thz3Wvv/ASF4ewzyiEiuKYZTur0s
7zp7sBt4xBuRok6kcM3/3N9Mt8RoNkwb4ZaVjVseqqEs5Wn6AilIYK8sRxdP0Xj85mpJtGRBJrQs
rT7qzgeprqRoLO4fopenzAw+DjqIljrZq2TyWgiTGJH3Po9xglDwkiGs0KorSg7EVyHJDPM2pjp0
hbk36Xv+vKYau0PajuceHj72U0I++67+1vY5ilaJaAdGkaj9up7kMZmoomylXlBxDclzO+5eIK0v
yhE8R7+LOV/0G6AIGaM//TU0U1Mshk7eHoSdy7h0XKfs6BjSaAJzijBvQzxIO3kgBjCEvHYwi5OI
78AnFASxzI8AeadqO5UPflHb9H06U7LbjlIzq0YRfcSakJXKdbWeOmV81wD2IU4kY3hg5TeNpBdc
3Efy6nVD8MJkycsGASe/kzcmjDYxrlnA6lcqhWT7istsUs4sNr7em34CZUKpwPuyjcMP8A66d9Vv
NuWPebeXnGMrTbIgUGnRnbGQ9IX+Lpn8whh1JrYqT6USDcLfaMdVEi3L9U2DIfSiRZQ/JZOj9H4I
N94ZzMl70RZSkiwV17p9XG0htKD2NG3pskhRt0DUyGW86nI0WJFJhz286e0WJ/0h8UNE9tIC6wvh
Fkgddp043jl3fHSKcax0mFez1P9niAAsddD+YCvlVnoKPXYSnlgbFuV5DTLT57UosaZ3I3Lkg+hv
PmsNpSJ7GlsZL6b9UoGlH3VonBejf2yZNCx0rvRPzUf1LHycYecogogBWGl64Gwa7sFmpb4bkNlE
mAlIkc19g2jzRcAYgzfZzNoMagrpyXF8pT+qnVPqgiq1uBNPTwlVg31KXcbtWxznHBgOiKNMWDeb
27uKcR827XxFmHakwmvG9QRLP+vzGFJWsllQbUTNPHiXqMwjrwxctLX1q/oL2clAZzKZCCO5+T5Y
fZaRlkbCbnEjPZWBjslW4kL1pqAny1mALFUmMPpJPLlfpHEc6SAcgCyhhY0k1awL2+fulmjFdqJE
Gp76VGOcVGuwrYatYC+072puwUVqI7yWj+4Ms5GhiJdjQ+ijb6W9qzB+oqGpoi390+IeHtFUGfBT
SM1BXapivJ4UXyKktZeMO3ZCJMobdxsgb4eXuXTOJk7DVSsiE9fH8b0vl49U3hbQ+/oaKWouCp86
jrEez/mTYe+KPyydhHeN3X/YBvG7CTfrm1ONQI6EyApz0QrAH8ipJxwhXbSThaCcaX+Dsm+UWFIa
IV46+1JN3vxghAU4CgyCsY3elTd2Bq9yvgsk1Bw577s2zUJK/j4NYhTE/DnyHdyVyKgkFPzEn6wJ
BUsPkExJyXpxqSfCzEbV5a6A6ii95x8U2VG1whmfb1WS9GCAmsIJhiEQpNOTGQAlns1YhgsBZSM/
y5YuafxoGwAZvE8aOlHB8FWkVz//SHmwu8vBYGuBx7o4AKl0VgHuzLW5ZCm++NPLFyH/8Hm/+uLk
QUS1r2CsveWad4HsMopYCsm28HIF+J6jmSTdKYFBz+d1iLwpa6NeWuZt9H05aqg9072ppl52NJ08
4FukSLymjUU/qB1lj4QsKTamTr8R75Q+0szoiOIFuR/DWd7mGCRxYoK5YsLEH4C4khGQdq+iXJyJ
wtY5g3hZk7E8epOkCElGMUrmho4JEA3uhpUREtigp6YWTVu2YbQ3ICcalOhF7ioP8NjrvXk2O5fY
h3kv6W3AbujHII/UG4J3H19DzwH6bvc1+EAlyA5oCGn705pYxXQF+bprz1D0WATR4cYnB2xhru9H
8pnAGDAQ9beZ90kvt0mM5nzvTMhu+OWe3WvPOPdm1cYYSHxUtFJx/hbE8gOr+A1mDrOq5O9lihnq
2rCWIgK38DbkVS2CWjSxsDssJk85aRHvwOage8FJAmNDXWD3YhiIiNIh9e8fvGvyzw1XfbifR2f+
/3T7bAcOzArwv/3tRelAhjd/CclisDqcSwFpVNDe+ouOhXZIsHIBFsB9o/MY05G9P3ksTRrVDYjp
HBeKIcJd7q2v3dQ/RkMSys8b0fgV1oGwSWRqfTshXRsVZZ38jaQ9Z33SnpCMjJd/PlOxOmpDHhVL
oRGbIgx5luWr9wmKYc07txdrhM2oxAUwc8j2Mufm35CFYn62KJGha4qg6f4XyyXowQeJy6lRqusl
RriOcowQ3H5l5BlDVbpyc612eQ8tKzUi5pCNPeDMDjOvRn9lOUhUQQ2+x64t8znarb3Qr1iFyedc
LaY71SThBRnArNDj+w9hft2DfMpakRjMxZwBNzThc7DM0/H0LBE8pFiCeZr7crYNeLisSiFguyYz
+kbbLPitKBeiV8bnMGGxkvwdfUnHQmGSkGgI4C2G9ejYUwPf3fR3ueVgQIGCAgP4FViv6ZirINYX
+5l6SmPh7FoLG90GCO5oVBjdOyOv7rSw7arYOxJWGTaxkV70qydLv6B7+VQEl/nd68uSL53Tv6xb
pTpiFF/HUTt3QB7FlhfwnohYXmSFO1ctT94qVuYhF3TDvucRQGvbuVn4+RFLJam5A1PdL4PU84CK
plFoEkYoH3Dw4hSeu55+vYu3qFyBkcGXMCGlfu++FRzo91t40wBFF9SXAV99YawsaOqY8LYyeIXf
7BwNedb3msTJN/ITBVc2HYBIBtLpmyUFAWXihTOqXx6SA+hyEOZUvSmxZnL5x2zy3nKMu7bEDz9A
nEzvRCC46cshxT+EIg9f0ZbflqZAdQQuSqXLP76UyproedAe9U0tZlUsjSMblI7uqPBa6Yugu32A
4WyVvrd1yfqY6X0JlCZs2vntUCnI73r32KOf/zjPPiKTiT7H0Yq1MscsjyAL8bduBUXi5tIGFqaG
mVuszDtHLspNCQ6mFof2dFQncznkxZHEhQzONt2hfCkSoxAdHLeezFPCPI8e67flRS/WMl3MUSTl
tcc8suVVa4cLw1+1Rf2vWJswEdI8yGl2zxkUGIA1UdXh6wXfJTZ8CRRHtsEtx269DPJ5zflL2izB
5QQFTIXh9GX0cXueTE9+ns/zkQ8lpXriZPQmiDMjJs/IN3JjlYov4PmKJbBcCOy65kCmRdfDwsRd
SBDL1h3hyaXFk0nJG2ltjOntctU9ETPDqBG5bpicos2vYDTUzbRoAwjZs0iTlts0I6Au3pwm7T+R
mcjH3YJg+7rGZYeZ0fNLJ/nR8LWss83p31+DggaGjuhKtKDDZCzvxZHR6etTxTSfQZ7zJ7ksDO9F
UsxYazGWC3SuYAduVkOc0agUP08reN1QuXebjb3KFFq9ZYLgG0FVJpv3DqgZJcjCIeldgdL/YN8b
Ij5d/PkoUEi6vw4qs5u+Kz9z6hDhDSoMfp1oNOqDrjKf3X2+B+uSTauFn+AcAln6ziNGKBwhqxcx
v+l+DQfnQP3N9B6V6Zj3QddvCc6bOZSugWRLiuoPdoVKBEVVX4tb2ZbioXpxsEi2yOAg2qsMBIxM
z5nGf0QLRswiKjnR3zU+hVQA93XKcMPWF9SMM8osunSQ1ieelg0bYibuWrcyzVy8vLYfhHFCUqjM
suyoTuiItvOTEzYUXfXYLD6kf80SKsfuo2cmsQ1QLbDjvJnjQxNB4rKicLRRocxrJKEbTBgltLih
1ztZToaXWT4aCqcbee+hYje9dZ2FqQ6iz5MXOn1Kpz88Gl/Eyi/aVkb1SPmC+QiKZ95IJnemrdF4
Uig8zjeJZv6Mc3Lk0YVOdBERQ7w2B7fl8D9/D6Bcogwo4+k1oGle01lgq1XCROkLEJnH8R4W0DqW
Xx1jjIJYJnnjsE16+xYs8xEAX6vHbRjyxWEJ9OB1Cng6HNY3hBnXhH4jnrjd3BKnpvnCB4wFv0bq
/6VH5xQ/KfComSA47//Q1SqZuv1AscvmKdLGEUHnAo3rbDKmmlZ6pLHr8xyBp4cVc9i0Xg/1NSUw
kMPgshtO8rHfQzmc9EzHUzaSUAnRd0TspmQ3pqSItxzm4We9qmq2LVMnPmjU1AjVY9Zwfpik3Iyq
q/aPEKDfuhdLF3RAOI8DPe5z57V+vt+rbI3avbEBV+yAu0Znm61w88dBoSPDIIiycvYw4vI/BvhS
8QgVK/xpS/B2tRGL/ENYGDvQXeqa7+cb7JOPOLu0PnU5WXUpToSDU/0EIy8v35VWns90a0nlBovw
je3cab76K6Y20RzZJLpGJN+OKFgHDVsKdmHja85ifrpIlv4SpUiZVUwDdLh3oJp5hQSspCnLZFP5
cQJ5rWIIkagvilY3Yape3kmXkB0z5iwjVkDIX4UmYCqnwGMYBsRUgeBxD8THpXDj4Y3ux/sD3Ju6
Yy3YBbfFZzxC73doHk8miQgCTGbbYp+99LX4kxol7S4yoLFvhrPzNuDGyLVJtL9lKsZCqbbpmZKe
0hy9hOSa1Fh57x9L56eNRMDSc0Is2p5EKiRLmhZOoW0XW0/tuE6EtAnw8SNy+rmYTTIF9zjpthJ8
aMD0F/eru626cEzItJ5EGiLEboYBjaz6vT+xbiQCfxSWCbfvCuBGPanguLWZhHFUBQE7XldwEqnG
o1ZCUeC+RB+K0U6LE1Khd/WQv00KqcDr66Ws5fLSISoV4hN2tAf37Og3jDbrLLMCOnNxVuO6UmtQ
JJYg3N9pK5+jDULEdKAFBOFK8ZiFl29MWF8PpG3PlZcmjWefMU7Bke4OuU6TR3B71EXLsc7YIAgY
zSP4VMOPaYHY69WXUM/bCYNB0/8g09VdQ6kxaVvYR/cHEQwsuaG3F4R3w65bxNfnsm9+X89rPXqm
fqs7+ZpJ8TO3MDU8hSfDFMkDKKR3Kxq6cRWALf23inKPX+Gnu/LJZ5T5jGr9ySLXoqt1kRXii95n
FLrCgsi/VQlf3Hx2n/BdCNc7fl0J8iiFN4iUSFwJ4DWB+s5VYABWouNPkTOYlwfHexrkgG6ALVs/
GyiSIQ8W0qTA7oxvn7hKCKiK5el5OOJNp67lr9dRlqZuyxP+R9tYUwNbvBC1XjUJFyerfTCkbS2h
fYCM7e7V7m08Z5d+0bZPu2Bc5mWFMQJdZFPT6yKlstRNglgCbQnIxah2RQhKdhFjhhQVS18gHvua
C4S/AO0ja0Ov24SA7OMoGziONxJXV4w0Jg0LfPBoDcWsEE7J0EXZ5E6oJR848iDcNE0r5pQwSIbr
xwOLCkKbtbBx0lgeeE9wcI2ZWI0hU4A9+4IbVMka2jwveMOxD1oG/VuN31RUY856It2YsE7AqmIs
XYyw6jirN2bVkLM84A1DtXvBzx9tUNcx2KKDznYY0uZ4tNnrWduSew7NP0175FYxt8EEjgFUglXR
0Mp385Iz93xaCuvms1S7Rk18B22jlsKELVqKCy1oH8drKbFbmfRPVNnsbgawgCoTmcethsF9EhEE
PWl4rdnM4p8al10+0BCP8sRnZLPWzNvf3pnTt/MfWoqvo2YEr7d77gASs63fO1rkF+8NfOZ5Acon
EZPLJIVB9Sg7HP2FyqqHpfpZeo32X273FkFHIC7DhIbWEC4psHlw46lEn8X6jncODXZ2M32XSuqE
pehJyRFco1zKVehjyNGliDFIrWOPbTpbhZbnYwgV+H6sVN7zRKjAoLAr/xnrdqOIXUS4QAJa9S81
DLBUKDvOVnKCGOWhnVDH3QOVmM1bppZX72+JrvZfVX+0A2ZS7sr0w4CXnWfY6ZUSzJnc5+dE+U4P
LXS0EjmVLnoxMjPo39FEdCRAot56OKAJeSXzMTEByaRI3H8u6/wcU2kAzp8UwW10rtAntjc4Kcjy
mzFNAEEwD+KNUTd+M7dLjqBwuM55lFgm5bvjQoSTjcclMCFXq7hoQy6h6KDVqmSi6nKU/Z+zL0ms
0GhGpXVJIPFm+VP2Le6bujreY3AH3jU902p17cgaH/VhyDxGCPs4kRfe9lA3Ck7dyuHJrojoyqyF
CPWy+jg3wfJUOCZHQf2vFlu8xEsW6mfMdb9rWw4Bz68Bm8ehm9A55pQ17Ys66R4go0LWgOmAAcuH
BVBfcu1AGzx/+LgQGki8D8UbiK8/5VkX2aBf2UMeOXkHbqrDoNdxExVIWYLmg3VdmzMPUTme374S
t21Nd2PIw5eVUDtacFSUHp9dgtgmMXUk/YwusAcaQG+wak+VH08L58FnjG5RKyX/8/i50faXq/oW
s5neE7dcAUpQ/5snJMm2dpmpucmStMTLbadOB3geRAxagVAXZrL7YH2Hg2nHWzNnIuie6PZg2Efp
hDxB1dzJZbBMiO2bK0A+WY/VDOuo10at0I5kXxJzE04y/LXfqcZFp5uzTxPzYfuFUdujSGhoUB2U
0cIhzxKI5FB3BxfVK5QgEVNlgfMA0UidfqB7GUqUssVU7EZpgGSieP+KwHAQjgt4qd7MVlgP89mw
uQ21YChAC3XSFmcFE8K2/IxOo8DoW/MsQAXobAJjQLaXymKk/CjfSE9JvBXlWaSKqn8FhByoMJT6
FbH7CSExrNkns+Bkw7rbP5tcut2hV2rB8E9QOgI0VdItvONvxeY5vOnY3LQ0CNWV7Qo/nxaINDQh
uk0gPB11Dj+PYKsck+7Huxao3q1kqlfZgVlFEepN2UvyGU4ZVV9d2ybcxsoJS40TnZomeMggNHae
gQb35X0apyk9+U7VIa/BZ0IeFvXBleAZWi3Sl9pQDKZ/PzD0iaifJucSwAGggjOubNZa3cInHfvM
efIPdkXiZHgqNaIvkEAkZHRKoUeAf7VXtq0jr+gUVH2qQ95E5r8oLiM/vLnbO3ZN+hTdDiFgoywu
trW5CbyGk+kcnAC6hZ1ovOS7n251gaAznDy9RM7Z+FOs6sIQpro7Sgmt8/ELDEwYqYSY93VpucRM
EFiO0MMkmCGN6q7sKzsgqPwGZb0UziT+211ag5MFgKDstgGseUsO0JMapegrOEtIQxrQFLiBvzW4
WvUUyt+ah2x5JxH6zvohVZxYoBkM93jG8LaeNBkZrcTX+tWSvCtLde9BS2qkeUP1ApbYKP7V8UN0
vlhY44j1sr0iRKg/o9Cu0gUx73jyinjcvnsl4nz81kq0IqMA2IMaZk89eJPSBwI6WmbTaWwwSrwu
JzEXatJNpQ77IB1eGJxk1mQ8tYohz4s2/oHVJtN8OfhfqLhM+l35CJmLO+J4aCeAr16NnM0B6IKa
xFMcbe/vCeuj1uqM6iwXN9MpYPQaHw5zmLYvOneZaTrkLJY08fM1/++L80wuEtH84NKQ0reFX8SS
STMJ0BOm5Rx/p4ZEKpjQYlTsAIlqeE4zAY69Qch4gdyjBjTA9JvyWEtn2ynySjrMIssFv9W1JZee
2SPnX9a+Gq/OzJ0dQH1A3BHYUnRIcbDDZvtTbn+wyVit8ye+8LZWciA7ws3T7JsiWux+ATsEOOUm
xY1G949i08gptsLWOC3NXhvGkmFmkfXq3h/9pR77cmk2zMcoEBLSrDQMJLzT8YVQ8+64P/yDevXP
n4XY+EjfafLl4/fMNI9v2tl0ika8G3TS8ZHbaQiEamhYRrmcJbsSrF6K46WkNefLVI3bK8h9d0eJ
eJN4psXOgTl3+HoheE60hjHl0M2YrmBmsAjby3srdPA/BfmcXv3MqzovTNQECngvyL/CcF818gtD
Kg5ccT6e9g2OzpiSPx2fBKZw3wn+H4puEDW9I464+mHHnUYJZB/I1hvzvkFjMxWEIhsa680RWk5q
5vWjQvj55f2MEIS44wMvtLExALz9E1OZ++gW7BE/wQbbXXZ8Kv3UP9P8chwy0u22Ux0nFXROd31V
kGLlCFeQQ9eRnVbFNYes3cmiJ8EJXSPc7jGIb72Frrd0gVO1Yyy5ox0HismnM588M+BI/hxrOkGn
fO2CmKI3RJE1g0l3ajRzC3nUyUiZDoNZfxtlLFimApE0BpAcF/bStOIz3NYKKsPO7LZHtm31Aqqa
arDErM8NJVv+uo8ovjq/b1cSWH20XVqFQFMrQxmAq1IhYfbxK/jgChEEYAjfFCuqWKLRa9f8zftd
3tChWrTmiAHmjuXtJgKTnolOyzPexmEqPJ4FMWo0keaZZJ544OPLg/d5P0dQAdE5KJhcJA1LM0YJ
ltSdVSSYpSjOD2jfjCzZ+u/jGsRChQ3ydKPBHk499fKmvJaXrF/rpfcIBF0FPLAF4OQTWR2fm6IG
ZKjA5YpnFSyulemx8TacGHJ0gkF7OWlHcts/yfVNvFXqcICa22CXc8CMjtFh3CrgeZ4XVIFGUVPh
QhCr+4H5FGQWzkGDoQQYUGzb8U2bMwCkiGk+eCY2SUg7VBay65sbXLsCYAz4LM6eimv/ldr1WZrz
W4nBeXnwKVdP/ej/cj12hShlw5D0YpiMF2f9CmG1FJFzq1cm4KGI9FhSeY97vPy6DF2QcdK+eI1L
bM/YcMScqcz37vtGHlxjbZ169J4K7DXmoqjn8IonQx2w0aAsoFNfEm24MoiRxVdJHE7iB4Wu8of6
f56Plpyx2akLNxJu/XFK4uyUT/zPpIouhdc9veLkPWjOI8mdUczplCNkScIP7UXwqDxNaNczG1wj
7Lm23rln7mptcPtOGRwwSAO52+PVdd37LRiBUWs9daaVQevKrk9HAY+OekrtqpqAn0ily3BtXUuw
m/vmDAkqa95UtQXm8Nk9ONQAWFfbJKT0fnd4QVwNgrXpxMaj7ifEFSyjmTLLEGmPlTLZeavSBDKD
aQ07U+mRQGDnmCOuOIv5xEMNRbOkkXJIMVfgf0pw9wM9v6As/dARARY7JXFxhdfKLB89QB4z7QW0
0p3PAzDOQhOjp4lqtVnOGTz6+sxXzUQTXZY6HjxcPFL0+KnYijDUK6lFAkE7lPuVlyBQRmZqBYcu
brjgD9swEBQ5PyTEz8RbNicLRcutNTTZq+JP2W07zfy8Dym+TFgS6CRX01GfgbCH4H+tkozMMaQw
ofoW8xIEdr3XNCoUf/VC9jfLHbbLCRJxRlnf33pfG+4upvDFe/hmcLxtRelI68kRIEauZH6beTYK
56o6sXQI+3d2z64YX5AoKys0hp3fwFVSmU41ZyO1gI1wW/g2lQskSOiOVj02AeCGMSObjva+1zfY
/TY2Sv3ySJgSxgG2WMBc3Gdu7NsQ8eWldOy7/nybeCwwCICw8PY18J9vskk6xNW7NiHCS3gml1nY
V4PVHHtu+3q82l0GnOptcVIgAaarbdFNbfMBfLAM1kCAk2kIHpQ5yCdXq4fdtIvbwx4765LsV69C
CIZa3VBCTgDTBssMSXcV1vdvVUvFCiaRBTegTMu7iEEmfBGbYyI9mdIHfqzK3Agvn2CE748qRd3X
xf/5V1UXmNFw32mw7iAuqJDDWH9ZKjTHLGIcjKA7BrZ4K//A0FFh/rZlX7ptxIJgno8RuHVGEpUV
muZYec1gaoXVaQTFj7GLoT6owCuv6QlxsYmVKypvlELcpe34UPXoEi5PgzF86S1ZiM6ZBF4qjiEa
d3+4c3QBjia8Ep1cdve3NukE5ndk+unic/oE79DWnvbAg4PrUC/ve1BWLOFfCqu6hGL6m4vOp7+9
yjY1ifW5hBrC9tdHLg50WY0mLVAxK42z7AgvCo4i7GNmMQneHs82NCeNcfQjr7sAHCRG0db/yqhQ
dShlRTvaSY8J2lX+v2M/tyUPkp4qheShmNR8HvoNo8TCNLR/oub3ovvs3JdVcnkN/kZaBAkp1fjK
gelQj+QQiRTGCrs4L8/jNx5cVVSBtbNGs0os0huJ3avWpRG9NGpj/PRvlgGoMYDiVd/WTTahJjyl
BzWEzTb3fRWxxUV1ST++sSFE5Fovoy0eGiz+8xKMiNkePePWsGbBUNwheU6q1qXQo7onOwfKld6U
8h1Gx/IFqNDiLV1kJPYJTKKSj0TE49+gih0SMGD28AvxSkVS27nrRX/z+vuS+LC6gR3yfXftFStO
aYGEUeVkfyQWBhArAAP7/PbJPkh9EScKZwrHfJcV2Pgf5nHOx1A0mzso1Ttdg8KbNsnNp7b/NARt
+T5leXdW0yEmX6fCaonUe5NMXd0jj0thUxWJVUxsHZjo6nM8/axY6JC4WJzG1Gv5k6Scs7g7vxOT
SKocyoAb6Pa4qzOq9dg1UQC4OmwvlQSc5XA8/s617wklia+O0tc90ZwG5yUJxSr41BG4BFYX8epm
N2LuCMu8jT6wSA5CbmnE22h5ntowOj5iJbzFpUE+OK9Wu6nNjUR09GVCWW4SGB6KoLlAu485E8c5
doVnBWdyLjOyCjGOUivTyiCMwtdyOVK0+1+lgzL4fH2ZUDnnZu548gP8d7JAVY1SP8GCYVPtmLfs
W0W6aJQH7CDou2CR5HZw3EVE/czdd+pW3I48NoTxY+/dnm0bWY9gahgoYQPCToW3ZxDhID3YGA/f
PqlcKn4QBoFoebsDm0ahK8iBdy3u/gB8x0ZiwMWFHigaJTPLD42pYuYBdHRgrKcu7+zsMWq1s/vN
DWrwniojbljCInUg2UUaGnFqT9pCthc9J/S3asgbdy6LR5Z0nlSjJ2k/42+fsDq0dN0LIBJTyHfO
TNeyeU49LspQ2YZ2ZzBFix0erQhFdYB+kdBd3OyGcf5qux39HBBrBNaFbKMArOXWM2QIiWSWXReK
p+c5x6NXkioCDlxTYxG8FBcdE3Nt0QwVO7t7xedohphF8ZUjs5Y3XPn5Q8HeVnbSqiM+WyedtFtW
hLHfHLVwODdLn+z5gaXXSM5DH8MGhQ9VU3Gl5Ao2CxOQPjyXT0bh1yTPJ2LJEcJjDSmaEx6ihgpE
kYhyAXEp1w4vq8ar43aGuWX9HBUWLiUOVBSDGNXhJrObhzaxQTZ2Iuq8nhMAvvOv+qb1+qZmT51r
tbRPeeHSOmV6bIP3jAZ2K469eynbw2uGX1vmbsjWk7KSkrB6Nw0OxL/mdqWgMH9T+zVhIQORTW7l
HXYO6g+i3c+yYMguVeG3aImJK0uZHdIpsDh/65yyJU1rAbL3f5QKSt9p3xv5VPIsqQICxcs7vWH0
XPZaDmROb4W6q4LPnTRHKnPChhbelt76A7cQHhrdH+2ZEBHKr0Cmf+75f0CWNK+ly5kMJs+leCgk
A8CSyHLEDUAXfe344K+U87ULYQ2x42+EgZjhqskrLn1K+CXF5MJYVl4WtrmOzvDvfFO1jKZpgs+N
5/FAEIezFbLT1fuAXBp5a0OGuCQ2BQNl7rAlp/ImuRvnixEg5BKRl+6eqvYYMu+k9lME74VqV5H4
mJE3h4J8fK/KwMqtIJ4+ALZiIGSoTOb7YIfDVGQA96BCsYA0jxv1NdOJnJcciG3AU2anzHArPYuq
7f2cc9/qDoU/phAXmmBPxEB0cRDPdBs6aCp4XGr3qqpSUw+fo6vVK8id6adRB7IfRoZc383YV0yp
YTybtkT00+E9EcGhIGTkOrX4R3kosXnKuliV0jHaJInUq2C4ZRLSpCkIrCt7gFA6izrhOO4qdQ0h
MNQXw+wpCMYQmxxU5iggfPPEzmwsOAPpolqm6hUpVm/r4CGhemT5ztL0lOewtZcjNQSQQCj/t2pg
BV49yavZtVIrJ3fzYNYVm52kszG47sv/71UO5GH/q7q0dRbwZ8AWo0Lp4WVROm4mTN11dmrDvJ6T
wysKLXgk5eVvBmU4iOwqM0ESy0xJyvezJKvDFyHIb5Ij9p1R61kKaaxCVFLokKsMniTRNyTvSB5X
YeHgV84ntCagjaw6ke9GI35sba89ntsGvI7Vww2dchDuWUJgtFSr/+m3gKlNvOfYE+CWquXwjd/u
ybW1WAKkP5KvysFjIjY+mavSsFYVL0j5lojWOr+v97iHzEDpB+BvhjcmBfDo5oxqiTMkHA8uWlaD
9zd4Dg8VYnvKbcsa7ik9vYMQFFW00ND4dnu/uiF7Z3QGSXoNxzaiCaxoSJ8xWpWBp2rq84L9K0dk
kP7J2BsAKWqPv2mDEdWNn2KWBMz7T9YbkezfsiyHHJDaaEcCoBBjsxx04REHHTd4oR81pLUwX6Hq
A2jtoc/T0/MG6h6h4oBME0jeKNREL+HNxP+pMaEYsYf7kMvwDIBf/0VwngLzfPMo02QK8mObjFk4
Jh998W71k/I60cvkIZfFCp1MgAFtDRYmPhyGChBQH/sYJdMFHUwuDmQFp9wlMYiJJ57DJbnrZqcQ
8vA2sUVtkK9bfX0QdYLykIvkteUhKrCN2Y35j3T9RgL5cNg8oAzhKwFu2zhRu75Ae33+N+lLSQBa
6BtH9usYgP4LY1jxi3UJU/gCLw9nMWvjDdQbnBZIO56ZKTpaQh4okteTqV40GWYFmI4lOuXO4Nm9
ylO+RHfYYfesc7qQVHYWhh6dOp6khlgA11lR/AzNFCpqfpHtWpwkt+tVTsZgc8DEIZXZkTs2W4qj
ugIr0GHDEhY8LwpC+IJT8uz6/GAeAuip/IBEIWSc9e+Vm5C8Q7dmlE4rSR7dZvGIr8RNPbH+DNTt
iZf8b8OzH8cYrn5nU0fXPjVvasPjWWsOboVsQAEaT1yNh61oxtJWwPfHNMioqomWu/VVwrKApC87
86VjTjsAdJtCjMlS29MQPoz0L8kBO+8wQJL/JGTgr5oAoYbxKQEXWODtUbWBNpHAPH6tUnd47Xz6
PxxEXaYnhAdEJbffTpWRXjDGjA/oQ96sviN7EIC712ZOvBIO6fbt2C5+QROeCZ9saiv+VWKZ9kgw
s1Vt2S5t0dEW+c9wtDZDr+d9FjdAoyi6ULT2sjZMUDfOvurlx2eCxXiA7OBVgvLgMniq9uH1ayeK
9pjKiChG8vp057Th/G4iPbqOlEkGWyAtnNQYPBSpkkvoOeIJWNpDBFi8QzjC8eyDWEkZiPAbZ4v4
nM/FYJ48mz2zQDpt7UGM+UVUzP3XyHtqQqdZYWr9+PsAOXC1qxHvlarWP5Jhlxn3PiIdfTRVR2HI
GkhCW0Q58S6VU+GfMWCZS0JvI0yaLEwtLQbWpq7eS2fOMTe2ZQeCBOQNML2QU/r3ZcY9PO5sBiDl
xidcHR/2yw51KFZl//aIJQSMPsMwh49B4TR7LBB5BBzddppQupmnJdwn6oqFamvD5nqS6WUu1rmS
9xPEyTZJ840b4+pI7Z4LC7SqNQuI3U16s+TDXUlaPC3WKNy/bKWNQrEFBvtBNG5W13oBoy/+COZt
A+tNZPxkQHoy7zyXfzDfR1DyCxqdnZzA+bm4DCRM3uruSczl3xFuLQfPL8W3fI2xV7nvxJMtwt/J
1VsYTCxoS7gFlqu5HqPJFo3mAaKAoHlxciaSv0Fk4N5Dd0kVE8ASfMPpZugnEgRpGPn6ImUThoae
HG9GsEmFjpxOWQXwTjc7GHIhpbkk939AqeSZ7n9ZxPWrzlTONE3RyUDk7jDmLZ4XeWsiZlKO3qzm
EdmuAQt1pKA2UJVxYaCoPZOrMOMhO1jYp+nnJExnHtFVuuTwJdLG+7Ns5SL5sUP5VE5ySixLkEIH
bHFlNODsaSjfkmbtatfsq6VW1BRe8fP/TLW4XPrTOlemW2lpWiGovvOL1tdMg2Ikt9C+gYV8yuBt
s8NCBli3Wm0Wc1uUZQ611zAZ2v1Hh2iMXpo7HNoUieZmvHTpkbbcTDVYpO4/EvTCEqW3mrzUSKpK
OEE2dxziRfvYfK61HK69UsmwwJkw6jwU51bXQUfJ+MHysBlWBvHh7sbxC0YX23MWkVIBjI2Q+YrV
orHYt3WNPRF8iyZbTb0WKLJf2vTN5TGN4Z4di516kQ1viEPRx9i0XDpbVycI4hmn6jT4DhLIw25K
/RJL1yzonzbW0oN7gihJXxOyHEZ8qQYRmBZWrzYhgJ7FQcIyt/Pa1pdZ1vu+vA0MLgGJkvNLhIep
kPUpa6eXuHxfHXveaR59d+BXMD4xsHX7kCa1qluElGljNUMKqfeN9+Dt8dRLlZms+i7fTZQRIpGu
ivI7bczxdiDXQofCR9B8dCStS5wfVSGdeob+8jFSUv3BPnLD8bmODjAN1qpb6ffcoRaXIGszoM2b
VblWwhloLer3PB8jLgtJqvMJxEzmn16SpoVuq3Mwh65qkYujlhMpGS/CYpDOPTBfOHNofQnDM4O1
/i70mtgOnGbZd0YHzI8KgCWgnZ8iLHy0aFTjZa1WeO4NzKSF0UWACsEkSdwSjhPjiApeEIrs2DV7
FNKGPWHnSLXCuyE/aU4nJZpwlmbsWQBfaaecG8l+TBzIWwY4uovqQErVwb1KTWG4oStOiqHJ0W3t
otjyiN6riRVmIhav3e43OSCZYTSUWavZauWH8pMa02iLW90TiP61CN2ptKIs2Illyk8VJ8NRQdtj
o28/GYtjgMs08IrwIix5UFv//YHqwt0ltWl72aMggcCllbou8xbt1Cgxlb92svM7OI+AhfmB25RQ
O8fJNc1nsCrXgfOEwOqr/EleC74O1IByj3sCkoe9gZsBua9xuTcWeZYcoTxS7KfsQgebeCR4cEKC
uthJYyuEGsVL3THjkTGQi0AvianG9c+mVo+Bd9AaJhLK/Yt4+WSrR8y6g032bzRfRRqhuLofrXLJ
83Lsd3EsLbrBoOd3xnsMHZojg9bbV7jbeRg9Ru18MT2B5Q4kqkRw4UKx+SNt2tQTgKQ2yp+llZA+
061NhijZtxlgcFL/5xCdtdCeNTn9IO8sAAYwocbQA14iUkr7pqQFagYujXaoCdaESaAt78yOZs80
xgEBhfVOf8dT/7ddui0jd2NPNJkXmsWNFzl71JdxvO/xxdV1DXWaBEcH3Pt20XvoAKkXqY+//DCT
Dk9i7NIyQr1isDE7DRxnwT+mOSKaCIF+g3ufAGVPd3PuoXN4kbsHxycGNdgkphaRE9SxQIihwER8
q2eppPi8ZsOj38OoBJXIZjm6R9wrAS5GG0eyskXjb9qYa08eYn7pqOvWplCsHAY1skppMOwgeltq
XCbHpjJNhuzx0iuSokT2uHR4Bt1v1o836WJj1ZmOeAVQlMlhuIUddM9dtqKqxzxy7vFt9+9ea5xm
azf90tvIdTgpegAgxUL04JrrpVLOmapQaAweejOVsqciGaInvGiubEe+e2eyDomHYSXRrYz5C4T+
ABVCSmCRRwZeqLpfVCg5NHaZ05/2knF00cAvdjVzPMiuMYXqhv0XfN+o+USsljO+5tUkPw6XMy8Y
GqisnpHacHngE+7AJ30TrJtDLpR+DJf3+pozk76TZhhVz2mjyP1f018E22qIgyi1rquiZsw7r79X
Ucb3mwwoE6hIl5i5ec+txbguk1jnMzPywJR53t6hrZP5EKgEPS1aPukHrvGEMK1UXhQqTp9P7/0k
6ZdonXZyUxZY45YRYEdCPvcNfYxBYOb/tjXKqEaDN8M2Hfl75fKppcYn9LpobQQ4Xcjo/YhA5tPD
9e2G1lKSIj0vb2H769Vtdwqg1M8iqq9iOuG/FaypKbMUrV+xeGSLjGZfKuFKK8vQQFQu83N799Tq
IxtPu8ABtGOnEn8QIZ0b9DRD59rZQh/SRpcSwRVsBwmR3fC8exxOoViGK2z8OXXyz9jSyAeN1ijA
lvtxGh5M1hs5wNRngQD+eyck7OAiHpbqgT0EcmwXT2Uu57RL9lnbm0+NI4oeUUzZWSAvf6CPUMVI
cLcBENBCyHePSAWKP0RWEvGYTKLXmElZwjtNaGktmnDh2NJP+7hKmIWSlKZt4pqoB5RAYemNoAfw
9E7Tp5h5GuFKvLerwKh4q6DytFkWUMCDK+/6atwhYp1bL3zf1gDc4yJVhScpGiJGVwI1Il8vgFt6
mchY/cSuUUfawkPc1MeJM9S5aUm8q9MrcMteUNXTm2azMt6SrH61+kXOhkjy3ZV3K3rgr2h4ZCXS
PVKNKO1lUZZmLaueK5URVHXtE/3KytJQ2vwvADt396+BpPLo7Xh3L4JFL57iDVxlJgU6C/idxxOs
EqIyrLSOSxJB44G4kL5krj9duNPJshg1yspjW3Cey5xYsWfi3KwUna4yA23c3WYC4VlLSE4gNkxz
72pkvnd+kinrjI8cSV3uDshbcRGif355hqIk8ehyqlLUKD2AyaefnYKUTGpAQQvCPX8x/Ve/XP+u
dsMR3+eIJgT4nv807UIbbbftFRKbXqrgKxhKGhULxUdosxwe6IbnQdkWIE1Ce052ags+l7HUAcZX
9Q5/jFW3GnjSKeP3w1tWLszeU74ZUPHkuN48oNxjZ3r7VNjsubC4NCnH1tVYDOJo3kRtg9tJL9rD
DW990P5sTrwSIPLpsKuaU29qeBgKS3qApw5wVFCjOVmWXcKkm14o0JBLv4XYogrxjxcoNIqbIAkh
lVKwRckQFwnMwmfRoXxSD8MaAWsWAzoQtJBAqGsQ0N6yCWiIkqNqvOwjpFCDuaYWuvjp+j63tP4n
kchkyiEHFtUuMnP526laWvAy198V8P2HMNhVHuuTYZ76Ps8PgBRx3dB58fSrx9IMnzbt7UFeTGrk
EkQutaEYhhyRieKYH6UTxB7jP7mHm29fRhltBdEFuo9EJ2pnxDgOYAEdFcjGT6h2FiGoBuN5jZkl
aDhtuNOTOQi4v6FYdaqDx3eldjaUnzhe4Xyw8gfPSt6dz6H7O1xD3f0Z7z4IuY8J4xWYmVbIv9sT
UhuYewrr3sBG/JAO5iCn6SMuZZtgQoXJrFZ2xqko0HwPXFyUu8Z9UDJkQRxA3tCLeQ9GfRn2tLxC
h0tdcK2N19FlFIm/+ng8lEp5sBDxOzOiVFLuO/MurtIJWSsFdGpqBkNFLkxgp9DkA+F2kFIKQ34a
tFVF7Hjhh9Wt++PLbxRy3//SNNynmJHI3oNY4eR0XHO4OpeTq0QUNiZVytErlm9W4gq/mmSlA3Pb
4vnL4LA5A2lsLCHkwjLP5t0R7vqgmM5iNOwvUddBiWDFOoNjYcPoUVoZrhnaba92y1Mg5Kz7d6WY
/Io+r+6qtWn3pmJx7q8dQ94kroo9mUQKzmbSZpLXMXKHFAKD2ZlazCLoFpBO40SGP/5yDwnfy1Og
yRfKJfObl3g3WCmRHg34fsAXeuFsUdpfzJaWnpTENtb2LVaLQ9+dDIcN6kapXbRtpaSbr13BJvNd
cbL6ZZsLDVR06kli9ATz8NXDAbd+Ek+vrV27P2LXIj0VAcnxQhkhdZm5S/DFQ8f0+MCXSbHGDBuw
xl4DfSPmt1xVufm77qyZSlnoFGsSIouYaaVRR+JQWikgpweXgUzY6TUvxl66Gxa6A73s2Ot/erNM
LqQl/DWwOR4SMedKuTNetB5TMbx0/C2g6bd5iaLltezpds710zGiq8KbLCDktKAWRiiJ+IWwFwp3
RkytdQ7P5GoZgja2686BYAKU9fUyN5KNjczMoZkLPIPKafaNyvb1P/i7JFk77S47Gx7JL33lMYpV
do5MQQroCdcUWVhFIpSR8gMByLPl1Ul65OttHxJdOLs3op/7sfLgPXm+vtT2FZ4h74IXOIAk1QGy
DQO7SDxCrb00tMOeEct1YtE/QAklX0o4i3CsKVOMdujpdW4wwIzBaBRoDut3jf+uMMOAPIsCiMB0
43dvovWJFSZhIecIq6//hJtvy8PrwByznudtDXZDCFTmjMUjxojRkOioO26jVEii/mt5or1eiGU3
0ew3nfnS6c1YuLLBEM6OKY5kduxaIbqWl49SRID37jw0XWtob0aAR/VetuHgBctXH2w0ycS8qRC4
9u3nyYPvuxFfjuZb+FY/XQD5tYIRGf43ovJ5oLOSgY3mxcxmanugwz0AQeLTPQerPPKlzOszSthS
AOsSrKVABq8Ismr9domkCC9n8j8Z25cclYeExKUm82g2R1K4829RdQMDWEKhth7nOQbfE72DzvWv
fahG2i4UYCA/jBMzpq4lYAhmVN0EKYGfkfl32aUQjuAp6LYC0m/jr0z2Wc3RFcF6m3Cr/EU+28QP
I9muqcdHvsbp87lubGdxvGI2tj8KPbrEGIXlBIm5xkKf0d5yrMpj3l/MoKriQQxjIG9XrrNVHeiU
NzNrnALYgmUg1wtc7BeZ2M+nqIdinjmufTMQ54u3oyu5QFg1AxYq8tOfcWMvtyVH+IJxWuTdxrHt
thKfjnDAluY5ucxgBj6wsI8ryKIKpMfS97rLfnnw9LCeKqu/LCfnLfFhd9SSmthC2OvqnUEzsHtZ
SoIzPm03XIjJNTUeT6c3Siqsa74Pvg5NasFSpTP4m9esxdrUbuuf5Wge5XCwiZ2XU7t+HWAqy/ef
9JsI1Ca1O1yOjaLUsW0h5xClUkapiZmu+GYvBc2j+AxtC0qe+vy4JXlKp4O+dxfIWEre2lnLaj9U
hSYvecWle3UUY/X7ytJziCMIlojoFCEOCpb2rfsLm1f21UPWpZYAONto88mRCimjYQRBVL1sviRD
POQluhgWOwmdniqRQq/g+tXJmor09r12lYaJ3xNfEa8eeNnvkC2PtUbKDLlPrSa5XLD6TMLjXrGN
p/0uE7zmHrnDupjBJ5HR15xgtJL4G168P1IoC9HRJd4rmY3dtwyE9FrmKnOtv2LKCUENMsgPR+fQ
MadKhln2sYpDpS5U0rnrLJLrgvZGbnUHsmfzFqz/JBzdmP7OrZeKIYSiZndoaN5kXEVqUpaleVIc
wdsr3NhTY97CbWBLOwQstg+k0NXPNa68Va+tbTHwqXu4+heujR2FzDlwte2r0V/tTE9gQVhUkaih
pBb5SEgXWTzp5ijVTg91fkb0IGyw0WnXb6XcdEq1dfxokeiY8tqZm2gM+r+gFc5povY17WeO99jS
4sn9FnuMzAVEAX+9kEFuEeDrYtaS7w82SBjpHIeR5LXpprjq0YXz0+5T7lDqdghRYrwZyjCoxyW/
F1ZQEouhcQ7Tn0/eD6h90G6VKKzjG6JdWeEMbmLwAyl4ic+bZaS4L48bbOH4mhAlulBhEUjAOKky
5Nht2JaWBW0Fr3cfKYdYLkpWvsxpuZl/F4+H9nSrb2AXMqzNVdrSM5ke1odXnrsZHtj5xninISGF
VBkkkGDrtPbQN8aYtPtOrdZGOS0eHrpke9JsBNHHZmICDB3nNxxrhJ8TS1gb+3l875bZqfmSukdD
l5g/9mdar1beg1zOVlQZa5owzec3VQJJ0FKT32yTwWlu90tzkno2tTBeb0QGrp7nGUpb7rQYLMup
6dC3GMv/9ObmaoQ6LXyKxS/dFQSsNGMnRYMmoB+mkB/uHrv2v67023/dF8fRWSL44jA78kwzy7+n
+f34vgocc/nMb3OaZ62klsnDzY0zmiDxzD9XiUXO4V50ZqKH4jZOHk8wuIrdNOJzsv64kISsp65O
2yRwTaxh3Tqa/FMb7UJXfekCz+02TAIu2c/u/Hmj//s3bipmUS6SyvKmMM/vWDayFJP+QrUDO09z
VIfhYErOrlAiSFvgMugCk35sNaNkAArkJrWtpzJUmzPgX+oNm4lLO6eGYt0DC6dEj7RTZXaMSAow
oIrhxyBN7FYBPlDoWUvq9gVr8KruYJhtt643PeJ6vnbjGUiEPKBt2qtWKh6bTtK4BkmmJsteA+8i
L3aHUUOK7LIUDxpwikddcUJ5YQ/FsmUY5Mv2S4k84Z3chyg71pqaLC3OujsYcz0oQjq8aPxb35CH
6XiDoNgTixstIw3Xwk8h6Dt45USe+f9pBx3JvByQ6zo2BDmO5jTWwFQTiO4ibgW7mPd75pbTI67+
0RmzuFvQm2CqshS7R2qqfDSRx2YeVIaaLPPcTXsXm0JvAwRy//OzKvGBcxC2y4ZCTd62QmNXto7I
dqh6gK93bBw3KfxlIcLALxjfZ6v8F3B+fxscFUCy+9VDFqTnJGViBeM/C3FGUybwqArAlrKRnCHe
SA04Ry+feZLxu2VyBAJuUuv93sngFfd1899YRDt3DCgPglFMREmvbCqBwRy5y0VV/2ECF3Y1mmjb
fKch/3Se/QI7PZkEVzuuuAOhBoBoyGvqfbqb1vLeNDVj+xCq+BQ6cya5dGytOPScIX8NoZTd7thU
T5XQNyF4S4UycxzQzOnjDSAlOrGlQ7PWIFWHhV6u/9hmdkTGorB8wzYQZOl5reJD9bWP89ZdpYB+
EwOOlNNqBKPvYFrioT4hDIAfJCET0Nars9AcCAWziHhnu5nS0KP0r8WQOe3wSjK7u+wOx+XQAtD7
lYShD4GIfuxpD3aDOp46fuDF/8gbncBrAynmWJtCx2ubSjMLha40zkpTaPMmBqt2wzFrwOgZ4lsj
bPrl38fMOH0F0JTzNF0nzicZY4gn/3vV2P82yrl4p3KHXfMyjsT0YKf9Uevb5RXVr0/M3Yx9zO08
jPTlmBDXZX0Dhg6mTM5NWWpKGRxSjTejuk+H6Bnk2yNlcmQ3X5zmGiZvfrENeO+FeP16XyO8zz4j
cpOFecXaeu+gprLf+GeCVYlrBZq+gcPMcLfSkXiYsB0y5blVwpC2veYzyJWtF1CfTxke87dWg1ap
wX6vX5j0OcbLYzqOixl7VWtR5W0Se1NW24qZvaW+FcN1xzUb/VCkufSQ527ILuCi+Klh+M5SzusS
WtZzs63aanlpSv02iiwxp+PL10kxJJ7XIzhWIY88fNbT4D5T9zH9JLVs/mqkFVuo1Ob14xcW/vOG
H9/UH9oYiFEyzINjqs/NNk4Zv5po+P8mIbnX8eg8cin6iaOSX8/XP5I44qf57AEV5E4uTbLvR+dE
qta0+pq3IM9NmPxAElT9NS3kCocGrqyKmR/pvpUR9jmDlH2AJ5Mv81w0r+YlGI6pT01HkjXZQ5S0
R4mTd8OuCdueZkwp/ra86LBcY+xigXGp3zLu4Tu+nYJ0gKohbUo9YSRZgtM8BgxAecBGBiMxdDpG
qqOOXwe1Z1jFAsf3KBV6H4RqYWYNcbqVqSDUkGHtgaSwpmTsNLZ7J7iZ4Ab8YyEZJv0Xh8EHqNe+
p97+5Y3mh/9YSSI/nYG/FvEqZzTvWkTVvX8qdnNSbIQvcDXu9U3MZci8NY0RwjS2zaqRzcktIajh
uONHnqpp54iDRyM0gx8WE6skEJ55oS/ccebg7m9HWryZKzfsKyLjlWGpohosjgA6+umqfmvv/opE
VbkgZpGjuRR9rOIBlvs6Ipp3y9riKpdmg3zmPzXAg0TRYSDuFTwEp25Dux35WndPzpYWeEzqZOvA
vAyCF/fLTVj3vuR+qJ4yAVH7ZxaFPygYTysV77IUfHhKvpDUxhsCawVpYSt7iMyD5T7hTjRClaai
hzoayevxdb3eEQ+H88RwQHU609lbRm6EamHW7g3opO57SkDZNVp+o5lMyUC7bjHQ1RVhE8oG6dFl
bX+jZuLbCp0rRuq2bNwa6zhn/bQ3Kx5g5lgrb5Ecq74lfmdmg+ESb+0EdStU9hnP4KdrvhR8GTC9
pkgn+c8ULkKF0FXVoRZoS2aizTvCKa0G4LEMhYg+FfNr6oCEQDdFwUUfOY1pzqur8JHgrRpOaI1g
82GAXRoYoGVSNcmbMq18SROyDu14KAM21naNUUHtbEfbKkdUwujkPaX96w1HHrO5NLf9MsxeUAOh
D+Nug0JKwAmD6Q8WkSk4XIknvotc3IBkgstyZ4netUynfUwQGzfX55xdyo3onZYhgOaJjqzs5kMt
sQCUER8nr8j7kIyBNQC44GUkuG8dIhx5A0AFDEVzodfi44lz9d+pmqy3YlRJbtYbfmF67wf2cr3b
WVB0U+OAv4v6WKIClEvZ0KSnI1LN/reBwRfwoKVz6uJPGN0lZxHLTfdhJsQSSIJTbxrS0YwecCwM
IlIITMUELoEp77e6nVXzGv7RofjJwn4zyOXCo8658Ew4qEJjf4LXALGemR/2TR8y6p+bYv3aeauH
U0itAPU8s2xUguriL3wrSkFr7O2jCSAj78LdqCI3HO9JPCWfgL2Oi51dhi3OCPPJ9YZeI1+jZvKa
HRp2D3HcWD2PB4hcP7zkujjCQjvoVZJySKTRGFwvS8Bj8JrM3Bj0t/RU1e4qNnPLpk70RCbaFKK0
HhV7XwYHqJIZFZ09eZv2wJq6GPrCE+pbITSKNSaxOG5PuiCg9+tVFqdMXMIVNpYwivs4GqE5J9xE
Nx6c6GqnKdfFsNND+PBCkGO9V5bksmUAGCY9nalvJfMPpEeFV2gP4H+mvItLxj4wp4Fq4Vry/WJ4
ku4LgB0LUNI4n07i3WQ6X5h7pwmEW8SCA3i1kvy/MIaomGbxo4mdEnxsMAWLe3rL0QMsW9/NOkly
0Ho4X1y4qAyHLAQeDkZCNNmnUkDtBeHVr8pPAgtjIlL3xFTL5QREa862Heh0fmEXn7rjbvLW7dvz
2yd3UXDzL2FVKRJO1sJqQsz/oC+8fM+MK9SqRWwjHWypP/yES9fNlWBqklWAUNQsZ4YH1sIyzKLc
ihXhFnMtmcn+liv0OPR32jsrcU7sxxWvFGk+Y2EVt+qc2r9QTo6WTfkT+vb/5byN82XCTOBBvZNr
GH2c1LcAg3XAuD/KVGGm3pZCkK5EETjnbArqBrJYjEftea9iTFeICjZfrpp12IUtOCj8JkdmV436
0VCb1uCVgXs6Q/6CdX7Xh+5mdleRiTfe8LG3v9oZxhfgqYPvBiRorUb9pdCpkzD5EHadlpU2GiK/
tPPH4uj+/9CAahjonBghK1qqp0sPGSe/3dLtzJTamtGETO/fOYZEKV6IrWexfmv3kGenC9HzMwmB
gpVvk6nIpfCy/wKNwNecFO6dYYoIZAEg71h4KeLz19z4VyR+j/D0t3qpaCa0d4/ZUWgeUgtILZKW
n7aQfHxsEbtMJTWRxBxZBA8daBk7KfKlyjM27SYMXvsTRtf10E2x5xLPmJaKK7UAnagVk3HZYfwM
tiYQ1kwtTDkaerR2PHgAnQFvjPtTkdOFwKXwlZ2GC44SNjvNrWNb90FWpZs0PRQLfZTs7ns1Rtbj
d+U7Q0DEQjUxOlA+ZlEQ2vbYBe4W+1cbu20cX8gPcA3biF3A2OMto/whwIBhW8dWM8/eT8NQfRHE
rC+jxBHGCLiajwl7hQgG2IHIla+3STO5LxBe8gtRLT3gB5eG58FbZ0qYKtDoGigKZTNeU7g9U5H3
Od1Py28WQcIUneVV0SuXabmOOKX7vPOIsaMRZ+bK0lK3vyvjmtDh9dpU4H9Tn/x1lg4ssGyYwxjR
1x1YgS599QGuMZqv/STmKvfxE2W+gXtfn1qobjNN04DzqCBgrzsgCeNVkPDG6bUqOaJWfnlDbrDu
gEV/SP/W7jmEJAem5J0Ad2rvaPztiqBeei7GbH2Iu8tkebbYabZbgVkoYFxww/eB0BoDO+y9aFQy
1RWRbPkAPLeVyojce4DV2Upgt2TbExh01F8crkplHmPVwd68DjIrJaNQnfyEsOWko5Cu0lVgcyOf
oihTCam8UtF89OqMOb6Jbo6NzvsJJj6AP6rjfYQ/0++30bi5fqdoyEk7ltqQ7YFhNAuxRqApqb2c
4P7IhXhu5U6TPNSKuVyjtiO4Ank4nzzwj9HGMYFDybzWqGuIYkQLigbjS+43h+Jsa3aFO9QS8qY8
+btXcndNd3KZDeDx/63qqCktsIA9KjKjWCVve/TnpG/wPYsTYy/V1FgNKD/QqnhiC6mcZ6JnJ6no
hszM+ZJK6Zz4zw4v74ObrTVlH4UDhHXn22XHAWgGrSyQtkFk7fnVCXExFemTQJsVsLlDtdNCqACz
Fcuu6BIWgatR0v2l6NWjMHkHWPEfmueyP+M61iDgDU84wHqR0S1t6IyfdqbZj7de4EGF+mvblW7w
KoTckJCRkPYZ/OOUhW4IhkrBQQ8T4QWbzilNnMouY4uWRzxoYTBJ6dZJ3FDH58Iv0Y7E5Ves9EnL
/o8A7uuzmGmRAcKvP2xSddW3TrsvfFsqPy6UMJy0VOf4iVKWXQE7w1gxbcazs04QkNByJfskOx2z
R/4Vgw7FZlsiHJrxJz9/ZvQiRIv7P0j+L8gTj1YcalBx5Omncm80OIEe2g86F/36f9MF2qTFm2gW
u1qIt4GSfjqIr+fi5t5CaQVwf7lvm+H/vvRhciAVa36Bsv8kwFsZUJb2eKwCJHl5w890aWeHoMbF
XiAtfmMbWSfhMp1E0vLzpokvb4gIyopv116TCt7VhW6Lau1chwlaN53BSr1ARJx9vBs3JA9UAuNF
/RJswoMohF+Ol1lmK05QWd+d8LhDS4vBbD39Wllb1Ygcoboh1jJf8awZdRTd//NqEI9gVbWzc1Fk
Gn+60M8X7i1oygchNOcNKefm/Ss/b1Br1aN44phlK3MqFYS5+axybXC3gQBYpidT+E19m6P2kXw9
F7IJNG3mVGqX1ZFt+K3cO7xWLvi10ZBJ2nLwDiydlrTMUBhmoGrqq8JtVbAbHpTQS41PMYk8Me6M
jny2H/p4RzacTNyIWopgktWo09fdm83bU5FZJPguf5P+GxxJS5SWyu/8mCjxKtTcCnD28OYdFIrF
L1utLZD5Q4tqjlHv4RFz1twYyRRDAhcVai+PV77FrigyR21QbGSwZKQW/21xlWxStRd7V+6lblkv
O6KFiMS9ldujBHv11PTQ0J1CoGWwoCq64JK23IWCVBMMpLIBSl3h4TyDaCOms1oR+ud8jOsWcFTl
KYNMk5m+O7ZgrRYLiWHOpFYJDmGJYdsarnQCiD5G2+1IP6gf66dYd01Wdjsw/agyaXwq5mLCKypl
hbdw/fL1tK5+W9qzyy/h4IrgTqXU+8UkKppifwVXK8dmsIwBy72OHOHBSHaPA5AaI0LilWk3PZwc
lN5xho1eA8l/p4Ofi2Aj/EqnaZhuScoSnrM/MReOk76d16JF8rvNBey/Ott/9tjKI5IIYCBSiWra
DDuW+hFdr3z3ETfvm8UBBe4EgLZvvkfa0I2Yy9W8qWJfM4z54mQE4t1iFX0kkfEvIbVZ3qAwKa8L
ya4OiXJfuXAW2RWQ+dqv3afk9GRkZgO9uBJZ4AedQ26IaToKKEYfDoAgCezuSz9TdoFsfhxaVXA+
jPdEAlxZszm/sYClKqaWQ8LMDK3iykDNrIsiLQQwx32OAkc+KbeOggLrczZrzDoJ07HnP9M3Y4u9
9MEYrkMHJpg3luvOa02VmY5DwQrGTN5E2lHI1uyD815km8uuVYurZu6kamk63zn70Le2JPaYK8+A
EQ3SlkCOO4tJnc+wrPfXkcr723ASvvBWw5S2gctmp+TUaZrlCPi7KlS6caNpm0t5WhKQ0iirDLWw
Q5W8/sDy5n7zkHb8R2P9tAImyVPJvAzkCm9wZuScEsKcODILtD1JIn2brEmAPTYSTmE89EP3zJXN
1NFA7tv6ukmWz1bCJ67Pp3dUSdZnrEmxWBqtrMkz71wuyJBm+z2smCTwvtc0XlgUpTQ1UdfkNKWO
tM3hKrK3LlptpgAVWOb1O8ZdGfKb5l8DjnqEvku5rEndiiTmJ+6tFnBOIB5DEZZLSO69UyI2olC0
WABVP494CJPtQnhE85yuW/vyQy5X1jfPx5hkoSHrhyY051XzmwEt2ltLXyxTkGtVWP+9RzcCZBDo
Bd4hqpNKaKRF4MBO6D1xaOfrCwJ60PVZL8mTP0fbmSiDdpkxKGShpFcV+X/Y83pm8U8Czeobcand
KWdSuQBT6S5uX8LBYssSzc9e8skTrCtHmhfV5PfclL+ECiysRaBqII29vJFO+477Lzs62JSuXKix
cIl6evgLwH2BtDdBHgGye28CkeXJGOue776kX11DTjmq/tl5AVaOOVNOI7HyF3FlaG/JQXRW4OdM
ZNN+Ow4S88boLMyvVqhVOpZhjALSv+IFPIMxuYlWh7FoFrtdvtRSb4tqqGAoP/175gCda2m+oOiG
HNFpE4TaX+L4ugElXGu9cswBq6a5hya69rpEhPOFbPPHf7nguuFqmie9WPSLlJ7xKQmnca1NGb4c
GpFtZudpM2Z67hmS6nC+FiiDRiZvBohKs9Lx9f8GJyRbob6ZzUoM5+LzUSIphxS6Or4CwC5YE1yB
lScsukPtNrCxU7tK1b+u4SVmdFf0TH0Rz8nDN7inD4IGa/zK7BKJLzxDS1fkfqVUkr7rnBmvDxHA
aipehHJIq4gEf1qzuyG1pYkWc+aLF9rz8C1GPYSmfdK849ndzFLbiW4hTWFcQ8vqk4bjXxR+s6gt
VAq9p0tFohz3xguP+nPH8wsUCM8X15j2bgDmvA3xPfrtblWJWJLzwwmvMVpmH/soXl5cXxptl9Ft
fkO8Qaxls3cE3W4xovRAjxmf08dSJxJGxq3yasVs4FS3VJ7c3xViuw9wf/IucOmyE/sW8GX7IxO4
Si12NF+BIkWhIrEbtgzodmpWMYJBuyYKy+neVvXTR4Zd538aUVQ9MFcrTVyv1OcpVG092OvDaaMa
72dvvKI2UamhWvo+eaMM1FowPi+2Y742D/4niuL+FvRE/zTQCm1uKcN5HLGxdoLGy6R2WC3OKJ9E
bZoW6AFBd3K2AMcrUJeKskLD0P8k1XPi9NGBquNHreicHKAgUlnxI3YP3PixnAikJP0LUMzkcN6e
IllhC3kMxZZLqTYgqRzCormY4pdytOT+tSvuaBAaQzMzDJkf/1Ut1sDS9LfwHLVl+MU9UlFLVbGM
M9jc+LcJMZxe4t75KYB9ge/yzOj8TfMbpmjeIgliDVmNRS6QL/g958MCrLaJ+UglmN2jnuimTNXp
VjuIg2Svc8Y49wkGUBNGUZBfKRBMocQ5Y+rRSHpJBZuXGEEz/d1wK0TosnIOgb1lz+hVbHpG+54g
1Rf5NGn+0QOcZsO3Z0z9WJ28tPZLhgGofSkX40vlhO/tH4xnOmmFDCNID7gOHL61T2sMLOLWFQ1p
JZYOAnDLp+BURKvKWp0xM0aXHbLaJRyc3GQKSYncDj4guNSDg3J0goj8VS/Fon47DjUW1dZC9XPu
HKnPBLY6slWtNnbktDtdGfptk6X2gPhLf6vr9VNJaL9XHscKC3PKJ7syBtslWcC28a3A9AI/WjB7
JZpj9o35c9lRC2J1M4dfK+r1eUK90YYFrUJEmPXNmQwUPtfLrmmw8NSDBbQLG1PPtOHnc/miFECX
rkqcWnreI/JhR7fEE7cAWT7Ak4oOhT+8PlzcK3EOpRAPqaSmhbHxP/Y84AyPaEfYHb3iOB4f0hHJ
usKfYOpRmiG8lh6vR9REgt3rnpAaiIS628tawh7jSmIhaefXcN+L6lFTet/ZfdY5QNGkD08/HS/s
oWEzbHC0f8T1X6xom4aI5pp05XUKLACJwTrkJp11GxZef+0QyikzIEWBEFNZxQvObJkQItFS1QWf
7dmRsUzGcQUiLyDtQ6BuJ52oCst3+HBcNd54oudjMx2ecp4sbAlzSVoz4Yg61QbehMiUl18qsK5D
MLTrMUiSXsfLf6Bm8vDbjrPW2mQ+luxh/Wzve6rCbbQ6y2Auda5Usm7zpqN6P1INx+bOBf0Crd+a
ASczRg8tP0QoLzzN43HBrjD2EBKYyHnGnOb+bbYktTCTYFS486LhZkbDnpxPWl1w9dvNdNXVd5MZ
YpCogZyOHqq3Ra3NgqU9jSOcSGDdIbPEU8UCopPsCyam45I/i0skux42Yxssxuf1ZYiWUC7dgNzO
kNflO2B2nmdE94Q2KAvrkxteqoOrLzIktmFtgO1G6Uvwd2q0Y35KYh+molQpWL04SyIU5UxE8jyM
z5pJH/rfNowJjCinIDk10rClPjCUuMVin2jghgv5Hc4nRdsD7N9zs0kHqXcGVvm8J3Xh7ZBAOA6Q
zUU4jGx/vFxK4rB47r9/1Gpe5FPQUdZ5dlK01I9AhXW03qPabMJ4h8GSHb/CF/o+bHfoFpM8tP3M
PziegHkpqoz8JlEOI+fDQ7+0crxblLHTcwCLA523xUed3Jc70qIxoagaTmzmY5wIaklEAfYYj07H
Q3uTNrEBexyyxHvUjg9aeohS6kky9t1xYfvQW1tmWBgfl2UVYAoG2WSUO5oB8IFfYQXFj5/uCCkW
ECr5pV8sYmL6ouy+TWHgeAnhpxO0aSMWxAqCAVLN+dwtFhmX+2eav8FEftXHoLllq9ydXV5lmX1i
3ltynuzn3F6/Q2Xk9f7X6CKejynZ5QtoRA/iVx+Hi88NFiG6EbFSCCyUsQlnlS5UsYHR4Vh2KCFx
dVTiYVMBG6vD/nxTCR776tjyoyI0Vl33PvPxlQ/ktdq6MvDCB4EBx9/0j1cEXwgSJ6r8XBCx2QK+
XORtqb01AI/FKlwieM1b+EP15TIKMuQl/7niZfRnm0xgMqM6i7ocF1ZgoazosZtOK+Z+uxxFBJAX
b5VAGMDm9+IsxuVQSvwk5SEY3tIBpTHMMpaHGspJTZVh7AHrAl2SEWMS8Z2T1l7iea7dxpIblzoD
bX2ognYBmKI1/mLeKNzElb+lCFS8a3E4WBi9nLCaJj/JWc+FkWSjYZcjkkDOfqxghXdSrCntS8mb
UiqhcXl1xannCzp/1YBu03XCtsOvxqxl4NHul/mszzRR4xaNhHwRLvjXaRURMpktzlpeHPAhuaX3
6Z6PJuDVBZEhaSuGikphRw06F10eDGJcLllKpzXRnSNV/HihLWsYI9jIWpaPHwKYtSGa8OIxBLct
Mvhhz504HfgB0FMp4fAhxJHGk4TRO1UGncVNxA6WTkY/HR1gvwcfFgo/CVeI+IBDe8omtipM4vd+
rB9Vg/iwdNY9eigN+ldQZz9WwQT+fmwEY8IMyGWni6y7OQAN+v0IyBJ25Gm9cF0EB4FhX1hkNVxy
MtDKTyD4ClGblcNxBCag2+fS9yiY++dMDGHx7E1Z45zP7t2VLljTcw3NFDiHOsvyCWuReJSh4aeX
/IGOa9jZWG0o7eUyZWK3MopFiT0wkGt/IU3hUUbFJA6+7cromlSvJ6nbk8lpZSvEsqOHAupUaV9U
d3Yv54OrdtRxIXtpMrFMbniUsPf6C4ZKtro5TFY5wkV/2ohJ9XiCtLOOUVZ5gocJcDiGrL/0SP2X
9fvx4INIxDV8pWLN2vkJbhEW7JB3IO1igcRwbB6izNP7TADEel0S6kYDaQnvSOOvZyAtxTe/jdW/
dlfusEvrdARf7nFMyTvxjtSLLNRFbkjNLzRRkHwxX5TtpRSl8MryAFk/tf7fP4TI9C3z7Bd8RgKg
XemgcZwoUHB+sTBwUk83jlC9uEBLMIgY0xfmc+uaKjnD0jJPmTOc2S1IB2Eef2erueYwDEaILwe4
95pqCmplZuAeOuCLnOYpv/gAgeGgW6awVcp7Eh6pD+pcAwBuhcBESI5ntYWwjYHE9gC1+OrYvPPZ
ELJ79N+3m/qrCoLvpFyPZr/gt+biUHck3uDQMpxl8T/Yk5Wj08NIF3k6/yAvcALNeir7pjne/cDu
9f+6kEmmNvlw8TaGCB1sxKrrD2Ha8lqkhkRyUrF2JJ8qg8RlaO6qBZWhJglqbg3XxJsUqdl66AML
hbSoM4n82IwfTt4bnq+gPoAYbZsWtEdwsoDW5faAT9W/AU8XW9IbL+ihR6VQIuDT26QnJqTLyeqn
d39w5DP7rkSxtIKiEc6vqDyG4aPBXFPp6oKD5W2wA4FYX85XP7oD6lrET1mWu7ncWT07BiC1J6ls
TejLyRnzi8h9U4JQyBAmd+OqogEGuXLj+jMkvlB9273VK86H+5XSbBb8YjddwFHkVCszCrmj4MIJ
Y/PWdNUvEBSn1/kmfdq0MD89ckDATleIQ98zsgxmyk7fi6aEr8gY2VDIg/CM6sqCfTi7wB6nTuKl
1VMI0UuaI+3+i3r6UDsMZ7/Ez/7WsVnKlfBDYqBszpuKWycF4h879WWC1DYOOsTiy5VYYoUkn7Dh
oARXigaLp2Ob+5Kk8clv5d+4WZKiF+bPb7Mty/aU11LJ+xAcYD0OdDjq62s7F6uu1IyR90gtzUpr
xIrFYUFs71r0GEsFrW6yGgHBBFHBumybUAPWUOHlfEfSksdUpV62a1jn0cXBGXTFB/1C66dbVDkX
xYTW/dfCt/wsw9RZAFkaCBUWIkvgTE9XC53NY9GtVg6mBZjKn6ZKBvTFVRlgz+7ofjSUEQlB3EB6
4Byc2cu/nZFOJJi34W8/yM4SwSGg5v2YrH959EI1PmmpQ5W1zwLs1UlN1fEouWgmoXtdhGzilN3g
AChWLCdl/RdMfhPiuApGypb9MrT+lvXPJf+yXnFaLnCMquhnv69redYgwvPraOiknyDXBnj2XEd0
PDGyxIGDS/RZqWlZLIFI9vqEbSPknspkJKYv48uh0Hk15g3o41mwcb9WIt1cYHWZtypZlYNEt2Ad
EXiwDocoyxpjBpuAlSQSyeB0/PO0MsOcz7UAZskKCyL7EbviJRO74a571j1NTYlB3yxXMs3g63EQ
7J7KNTwsozZyb6NNZ1qJ/PnHjiCKZSbeZYDQVg7j/IGAVkEbB80MjyaTlnemeTdaZjwCc2M0vnn4
EVaAteE33IxfI2EB1lV0lUJfCoyZ3yREQdNt+CD8fchOTB0TMqz8QziM7h8VfU0zjwJ51HXOWIDo
XlevVkSQOeAHVE9EXY76RhiBhDWKvcyml4BA6Yy16622QDGpU8AuIwpSl7JWeOApvsiGRfYf3/UD
7GRR5M82BNcJGpXg8A0voG3VPFQs8a63I4oSvWm1b0Sa3QTUM5FmsrOx0Pc6Dujz5OfJ3HzqbxSB
iXl92F6dgU2jmxgXotC3oYLw6G+w/GrXtM+AII5biqy3tJ/GUUIG2G9d1FrWHuHForMnWbMftLCV
6WIdzXP+yaSc+6mMqr62vGjCQ5cZuC2f4Rv/QYnaunC8SjoD6njLJ0TyqrfE0ELNv+4TzxTV0YlR
JT0mvjfir0Ei+tQgWD/yLpT4G1pM0JTFcj9AC/YcsHPOocL/0JXcZEYKl+rCnMa48NKSkd8VFism
shJ5Pbht3u6IEQfGQCi4fZGjoEskJfcXtLdgV3eRc6aAZOqXL9KjJ/PcEeUOI4xtHhKOJVus25i4
kznm1KGMPb8Lh/ZG18u5UdaVHkuy3Lx6DmMhVmOV+SJgG3E5OOFiDp8WMV2EHXiItzKpyYfH1suu
hYAdScBWCZmvGyvbvE9OANpNuSkH0cfBqjhH5GAUyXUjguwF+iFvjiuFqBEr1nz9lTmnTIuVaYax
u/36jszMd7xd46WPXE8K3bK8scRFUiUBPLM08QLmCXpPlN7epbfLeCqASiklWx/R/Vm/9WWIYVtc
gvnA0cMajpy9n6y7IfpJGIbgN9F3yC0K44ZXnQMIY9JMTvDVVgH7YlTOiSQHQuRT9DcnmRv7BHxB
56lAVR15jH5QPHNF1egyydsazYicfAs86jfg/LiiGh7ReHxr9xdGl3fFReoAgOlDiFe32hCyrbjS
2G76asKvvpf0RW/B403QYoRk8W3MrAN1nZZVn4q8vRv/v3ckNc4G1BRBS3n04wrrxyp22F64TmT+
t+br48R5B0KDxLJJ1RK2GR02ik6W+pa4EV2gx+dv6wPphpPXZcdDMf/Vf+ccxuvI/xvd3s48KGRN
ldMe3fXs1B+xD/+9ku7kHKhTBjnW9LPsxgjh64WURZ0L/JVX0/a2tHGAe9aK6Z+s62tApNmoZ6Pn
i/5aBD3LXi7hoGAgrvw9Nvs1SMi3F78t0gXa6xhYtjigUW81sJWwkXMvWQFLA2/ryidf8dzFfJpO
luT4M41X4ySm/qzKT+FJC72frZqyd6M+1109Pyc+bhhccNSa7E/De6Da9bZLiMyHvkVBx2FKWbzd
fzCfxGtVo/Y2MqefTnlzdOOWG9RPqqtHnrSBz0dN73u1pi4oyTMlYK4kLrnMhgM0pgmo5tFC10w5
l6qFtEA9ZGaYeghiSdUqXclf9RDQA8SLI82Bv8Ua4qOymOXXuWiDjvPn13za9H4ch9EgKHNe0iam
ITNkzY15uny9gag1aFEb9grhDMUvvXVraZBmPAcZ7L1An0ViJ0seF+tMrr1qyLR3p/F0YS8bHviM
p3ihcVAXqND3Y1ZCg224aEIXkgdpQzRt62i6q+nsb1e1hGgbBGYH1pSTGjfDdNKHBT1yTjwNI3rp
jcazW/0A+PrxfFBU8lK0cK3yn1bYXcnCInDLdfuSxJKhKjTKJkcHJcq5ulefr3aKUvRtx3VcRC1w
wHdF9ZjQ3vW2vupzdW3+JUrdDxSgBBJ/rVQ9xGA9krYr1jQbwA1MS4ZgusswXCbtNieiYiKqoadv
c3G5GlQvhMzfjw7BdC+SC32fqrTHARdK+2IuuW6z54XWhmgmLd/dndjbhNR5P+ot3i10MAqaEYMw
uM2uE3AQijfUIy5j7ouGWLE0QW76CPJHaT+c4q/1kIitGkBf8v77Cwaz5aBcgG/yG8hXKFm6akPI
/Xa0rhhoy4okZs8fR0x5YXNvoE+41MCImfcaNkuuC4PryI1z5Khgke21R7S1P1NA/sk8MmX+8SiB
W63RMX2kxlWIeHeesFPb+hv3EVIR+iIdGwbSJwuB9/Ni8C+aP2wEqruAsaC2Dul+02Rr0IVzrM6c
gCgf8NvVG89qm7vmJEsMsyJFSOmtIsjbNbry9j6QaUdwZ6OGTaJEamikdFxtP/xsQG+ZgRkVERAI
eA/yZvuYncRoo/bVV9nVmFPYXNJijbU7I5Mx1CIiI2X8yYlrTrEwOnWjDVExRc56wR6lasVa2u/G
noG+LeA3CRmkb9fqWfNI6mPl0jTah5dcZgcjSbAAF7I+fstk5k1KPJe2HkVCt+G8mfJVrmHT3fPO
2iKN7ARJebPYMElXCFZmDlZ37wfSPkoWTTurn/pSHL95nYFDqpQMfLqA7A5t9HjO8hvvrJz17shE
QReQk5OuF+peYTYCah5DDH1fcHiyrL5gvUv6FOnhpZh4ss7WhfnaSW1qyfx8dUxPOIU1a21FM40N
n/JbifXKrOe8/Xc3LWnZU1rijP9CnJYWKSSibQ9g3baz/B9mcY1LkfEGZpA+j3vZgdic2nmC8zLM
MoBJW/bIwpvm5kWsNTeS2V7n7cPkb++8s83Ej+rVcFFNcA7C0lrJWXFpKe3OEOB1d8tI2BuM6/FR
JLgRbqCjNK4+Ahto0aHe4GAG0/NxeJJvVy45/hMQULnAfEQ0XBNztaCDMRRjGG+l/0cfUvn01psc
tFJRsc1kwAp62QQONBlQrOre1MY1rK/RHbwIWilpc4hdKCb234NjcT+q9tC7PxEiH2RY4/126CIy
iQLxv2tqP4723nqQLTMfjfDasS/MLnwSd3AS0bCiQQABg//XB//iSRGZuhI8kWWxWPpQlcblWqb2
CHDqheix8mwfAViw7TEE8UoF0pFsMgDflfV+8bD3zlrnAnJ+KlhQ/Qj8WVfWGV0u+/3UXWkMQ0I5
IVFTI4X+wJirKYZhZ+HX2Sfx6gtWpypI2XqEOotdO534fbMNuAax481enuIwDQfFNJ5bO00Zqlsm
pB6SeEx7kFKxcwkJI10etkwXzIiCWZcYaptHazMJaGKXRG0FIIpF4N1gXFi7WN/CbEbwTgWrePUD
BD7vdZM7mlszvqt/igpL7xQ9EKel3X9OKcmrqgq4ytl5sbh+Q1CtsKxUKmRYEapeWGt6jA/gwWVI
bcFgMn7R/NmGok7MObkOvclHM8YaHp1ChAOFxwF9pD+3SCcwyNjnr0GoaoRdoQtbEKdFOqbbx+Yq
ZiX19i7XsgpRBT+R9R8V+3dIZGimJKWMkaGCHpLAZQjn9lKnWvgnbi1xhQ7vNvitr7buxzHu5aq/
0RKya6OhuyD/zq/VQT5XAmePt0TKxK+Qppr9alnlXxtnLTAImb11iRZiTGCkg9s0sI70VESFkFC8
75ApbzOytbrX/Lmu8vN2rFnHorp3CDI1XPV5qu72DBZ+KedIab73D23Sys+1axEKcNyfoUaiLRNb
RwR1cboRMRRTqhd8bEKabNwi5kKKjSg3YiK2R+MnfcK0/SouRgbsraqoHN0267+IboFYfdABw662
IMGj7LFD1svjgnX+oMXECUjZSouTfoaQNF8FtwOENHnz0/wZHqhdLoblkledSMsQleTTZj8501hG
0+HOoF+3AjBhqaGkjBvVJpIb0oO1ESZfyB5tndC6epg9PsvnMVxtcIk9SOooN5P2neBjo0Mdq5YG
8Upvepeb2W+6NnRbEYwOgChr5AWxga5e7AQFGnerAfGXDiVAsCJy2f0Go6H/TlIh/RbHaCTDxwun
lUrf982ASvv8fRKhXZDeH0ZjHC0q0qTqMN2LJfYpqAA7eDln2Tq+u/PP3AeOWTQbrfiYnVi/NNK8
JS4KNq2Le0ZQ7gwt3ASy4WryqAsCxudPhgDFYvitdqstHZj3PIIiNGfRKW7QdcX2AQsyCQMcyOOG
eOO9qPnRDEmDO890KrO2HdtP1Sb0pOYv6Dm7DVdDiUtA/E9RQNjpPQefBkrXBunwTvZgdbm7FW5g
5eX+gWkyOTuUL4fQGmepheYe5EBEahLIaEeIBGXsfQYV7Jayg4ajf6Ib4pl4/4FeF2mepvlgS63q
DucQpwYLtmDxRj5m3yRs1WDD7cSOOFH1RLgToW+/QflMJJwpFWdKaFrJdULG7kt9ksE6rDSeSsMm
gd/ac07PtNES3uYzlQgBS5qw8R60GrD2dYYZmXsTAgfhvYuUSN4e/ck+BKXNuTRuKKnluiTRYtwm
2dsrJqajtpDX4lMp3OM1OLpqA19OBvtr920RI0VQATdy4sDGrq4FVWkffYA75dzLosxh4xraC077
FGGiU2fkN2lZO8SdA2JEad7ql37bvJkwNDkrAoSy0FSSV9/s2+DDXU3ivlXzGq+nQSH4Zsjo5Wxt
ooC+Kw8nNXVxt5emp4o4HEgv2as2IoGSj/HGEeW1ZFZybfec6aichu9SErQXsLw4Mw9UMYgI/aX3
8nIpa2N3DncTqn+MP8qifOqNixHYPMrZAl09w2iI+ujAbx6khBgZUWbskSMxpkFeQerebhBUdT3i
G37zrThLazMU664gKS9H06skuxvrmPYzR7NqZiTHk9PAbbIO/CIOCiU9wmDAUn7+94IIQf8Umasr
4ynb+qLfBhe5U+K0Mcs/tnY9iiX33vVExhsMXg9VIb23IMqRZvsmlfxwOO7kMJoqBZdZRxUWzNWO
8nJk9gbOWtleP3PdS6DR3vljWPg7fpMVsphF0v7ZyCXALCLxIZi3JcQdWOJRAQCSq0ZpO4TfWeQA
LYux4CWNinJdtEMoZSOk7MmW54+eyvNIFKHGrEykE1p2Xp5a6KpUAb0IRjPaoe5eEYn1P00Eb2+s
xtHOWEe18hcp9hRA2VlzN2DI1VhtTU7PcNaNCReHoz0zxph5JQnFx68DW6+eeE76J4C+e2G9OTI+
eSGR7eS8/KKdL/39v6rRloPuFoQ09HmlbZD3Db+HMcYcmFGdDBpf2MngE9Axw0kwp4XTHCL/3bzP
7XLvyGfXUwjNAIerOUy4+v8lYwXHI+lLpGSThXrJNJJluxjwkBwyD3Df0YcOgppkB0QtRuaKWoTO
7is9z33oPSlfI5XbtF5KLOzv0rDPPBF8HW9/baPdeozkps27cSyjynr9rAURkqdE27cLiObFSMZA
WG0g6lgVofe6+vEtJCGwazL2myMfKZVdeCN521jQOGCpTTS2Ztn//+h9zUZR4IxPKkxkzQZVdOM8
fF6gszscRsQhOXDos9IKJ0irzDDq2uW1UkI+d0+CbJ02skeUcO6b9HduEGtDssmmG8Sh68d5PvvQ
uj162PSS+BO5mLe/Q4nvmdtrwRpXUkPJaIwsOBGxOfBtWM7zeV32akxPEJ5QxIwGHchySKzVk66p
laqk/ARSr7oUFYtGGzkF8z0fV7zs7o6wyeLef4futMavasIzK+h8nnevuchFoSYja7H1MudRURh2
CiF5Apf5FyrIir0o7EC6wqwPKuVyDZBdG1o8pj5DPe9rVfzO8Px/kT7V1L/SfUziD5dp3764mO98
XHQuhFNf3ZjE0IgakCoh7ao0bNa5sRcmKVKM0A59mEzvC23Auxn1uHcGU+yWiURT13Hlgb16Qxj9
U4IpqAmrrLGBY3hi2C2Q3D18Fp6ISKEEkP8JYWZTsf7iu8Iy45+aTr9GksXUUPjt0JoCwchi+nrh
U++SPYDyaJpw/KZNfR84jmyT4RDMaMWkWrIRc+epTIKKjg5A8KtBOXYxRyZqhZCNksPkJ2jGhsZA
DDEzYOG6BWMaGD3LVm/GpceWHgYKkBOkfX3ujieLWC+/KtENs8YasdLH6kI/MR51HunHFaIZ7+6G
pKLt8AzF46TzmikVdcpFtbIQWkL9IZw4QDlq0y1Am1vIhDMTB4xZnJ2gdaEev1fKhm1T4bPPvVZZ
I1AeiOQ96VAtfzgUR8H3bnCWVDMmATZGi59gRO0U15vWjL2IZFoSytCzwtjRu7pWMMMN87cmK+Dq
I9t0h80NNeQvRqy9Rb8sabPW5+4lTtnFB444frEBnmh2wtz7TKvrI9JJ9OTS/WiE+9P0eUoJqQq/
5nj4gXZKYJfVx/LHRV5qPkYm+hwfL+kLT/D27loFE7tJpzoVzYxkHCTBuap7sVPdSdYaE3HzNqgu
B2OK+ikX3E666D+xwoYU/Nkk7uqtwvHquk8DwX7q0KnkFOjmqMFQYVx3H/GpKF54oP01dQ/GeQmi
5ErJSXmZcByQ+oNI+ok6sOl7RZHY3VBJXGI71/ARVpYmj4a2vXWDtx/w5q59AgNgsG/EDZJAEA45
BvVMZjRNzGL+4N1+oSuIWZvxI7FGLhw+faZ171XBNJ/le4qe3UFaXor91rqlKft+OCvwCHeXAQcE
J+5QmMwLpjsSSW/YeklWuwlTtLjS0l5r0wOxdGUbvzsS6dX+3VKxQFZQeMTpUSejL/AIVl8YXyR0
Hx8XhqRD5KfvxnLfRApyltklFcwMAQwl1ZDKJZJz3m17x0jv4Gdjag0UkvvA7BfbiuRSSyjzfzKJ
QC7vE4uBJwskd0WyDMzqsHB3om8S58eTvXPLXbu+ZQEoaN1wZCRJIaXVgqED6/i8fK+ARRYThfdW
NmzBmXh00PstGCf5kelYfiautGC/xj/6Qxu2kTaVCSWR0wWv2KHuWxD6tVB+iJzbphQX+2KrmJfD
IsrdR99jM2OWokDFrNR9ZgkgZnRd8BMNg4i4uhCkdUTdiixvK6Cidg+oq3+1ciSybVq8xMmX7XR4
DT6Nry9bksA9hEVPErLfmFLbyVzYM4Djq78T6rzc/tQQVhG12QTASetNGvM8cERTirgyjam85tyP
FlBBQUm0BYjm0RjoSHDpCkHVjZv5eHVGhdQhidVKkRmkI+nXpxzAa2Y2JJ+CxMhQ5M/EkK4dpSfe
Uvzzy+8sjH/Oxq5uB0Mfo9U84LSDbLszrbpOHnuFM8rDTspMsFr7+Gg/L+2Wlcd2vno/sBe9dB+i
PTbjQ354pZXZmn1pq8yK1jJgDu0QJaC5q1v3Wu269EYaO9RzUrQKjoZIkGK0ehKkyFZl1CP4WPcy
0O9cHL04sYgCRUk4ZuyahT3ojyhIcyEDCbKxYf1ItSBCDdW7MbwtDzHCms0euhrs9rCFLUWkfbQM
CLNnIrdCjACB5UKyi96/p+N8uHHUa0pKgjBWP1fN+lem3lkS7Mf3htliQT/S4tudCmsunhxzavnV
wrbkqcVpv2KUT4+pN6xGwqpoRisSdp7JCiG+Z/msvMYbjyxey7d5fX636bfvoaMPH6P5PoHhJG2/
9NAYTdcqVBmFp2VETeg22kvzKbrzFO1+iyyWmaRS3Ll8tbOY2/FfjB6lUoSO62PZe1cmyKmuQG26
hpWqdfhM7QaX4jacoc+cONsGOsLbloaArJCSc2L2GdFj19OpYWc2dR19bx0eJh4IEEWJEWmqcsna
+fDMo8ppzLrP0x2renPm+WQlhZTssbgKI4EPGxf4bLmHOqhmXV3SCx3z8/vVkUdOjguKq33FzDcm
HpY7cInUEAQ378gt8GoiA5s7whFJ2hpGf1Ns/z/uS5zveQgV1K55qK16IEbRPPiwVJaWfE2sHWB8
pGV7EA0SobxCz2d9a3bXT/RNIDOq48TPqAf4b0vPLZAeNExDNGHCnp3e+MCK6h7Di+k2DzcUg4lg
wbq4NMHpC/AFyCFOWsq2HiB8eropdn9KsBwK4ZIbuUeWBFdkUjsLac3YN+Z/SDpud/na/0kZ3k21
McUzT0rb8Yel5D3OYXHuLGU2QIDiZq2C2tncIt4eFmPF2iG6Si7VJzqILzjccgSB56I4klh5wkMJ
9N70/xpJ2TnLuYrzAlivXKCV48GpR32p+hVD6l1KppyJrGhUPmrCkkaiSdNqsXrIqdYMduxv1Djk
2/jmF+DpmlgTGZzOlxqGgxtvtwqyJgXit5H7xPJiTS9CJ8+AmxL1TZh8SGCQZUtfTsbsJgj0uwfX
w1S9VhkRK3wYU9G/7W27LkF19k+LLbhSCZB8qZocQ8P/z/XdSn275DT+il5OdoZrYeZ01kIPGicG
GUE/XCRsKK9KKp0ZSOWg1TkUtk2+ltTxwreUCKROC7dVMamgQWC2aQC/V5vQJQXizFY2qskFgMNS
hCoelNkEM+v1HNyWL99qKcEiJ78vQ5zQYiD2wapxwWFGHPnpxPgs22ns/Af+tSZteIjKJpXFQCN2
FnREZe0IJUAAsmSN53DkZnQEAj3hVx9jV3Cs4JucWa5rsl+TUA5BcWWFIHNPLxdHhViywE5lyJLh
mTVjWdO6sIKnqaZ8DpRXSx+H0fxhDBdLA+YeQZ/sgBoMQk5sttWVCpTX81/MgGK/cKBDNwgCWpvP
A5xjlzpZCDh+lr4j0GHupf+zf7izhpJEfQdFAFGYQMdvhfj/KNEpUgkVkDXWs2XPsnn+tyAC/Kbf
3etIumlG1ikq7QiP7stRfb+TaOGKpNNToftl0mSHiIF8z2GhKeBbpS8773afyIAxJOnEM/YF6LU1
FD2/63ozokjXZqAjVOjVBjgialOqCQXTMzUUqI8f/CGIM0xPgQVEq2dMREzLgj3O32tlnBC0Cu+/
Xim1eqeJJgJNZdJSpByBnZVfTmyxEW6rzsrzqQ5DCB/nwLym5oRAZuJIllg8fieq7kxOKZLm9vpR
qcrxiK2yvp4VsUSO1NVe4gHeiht8a0SQjcx05l1ogkO/9XX5w7UxDpPTStedo3Zr92glkdNPcRHW
O69R/5GGK6Un4tuTbzAHReqoPnGQaH7d0MsZrVeGVBSgBCZs+xKPBdARNjiqhVsFL3045ZeAvKjt
mlGYhGlFaUWL2T31CGopa8Sd2hGx7EbJRfJbHRMOPmXCv+rtdmgENe8JCt8mwSx5+HJTZQzS2Q9F
G3imw5YiWAN3pwr8UAWwrcT1jAsQLd3rl+1bXkfKEXqruiICMll0o7ylJhb8rdv7WwQg7CAvpZaY
wyF340wZMYUEdVvFgOPQTYaHsHylHF7W1yORgxl429mTHQpobSY8IYVnFTi2/epd10yj8w+UEHTd
Bj4pfPA1KJjbSHwDZ/OLzFV8SL4XG15UUOx9PWii7E87Xdw8fe2XgmX4eZdkyMQxpP+Kw62IpK9U
qmG8rrPsig0rFIQa5P+ZykNjWWbeBAau7m2vLGpS/8c5mw9KXRugzNyi7tdr5BKSjY7DF794fez+
jqcdbiqWqqV4rqH7f6U1U1XEPCj483tAXS026vL891aCUME7n3tnHFp5juhT7ANPZfa+OW7etZiq
QnUWJ59CES1jzce2nZDrEPRFR4OWTw7aF83Ig1JDjQ3pFa3G1ULZv7VPLVhnY6r5XEMX3Ccb6Emf
wbNXCf3+sKKj+Z9RPPUDW7uEb70JnDiKR4v+3Fv5mO+IGRpk/UthZ+UbUPyvNSW1pGMcxPkMEZWr
lMlZ6F8R8yHX8WEZy7F5k48FF3Ws5jtuHZkGYhqJCOkv5+vJR9A0Y3C/13ojIfEWq2rd7x5ySPMh
OFD47vQxW0GumvgVSM+tRYvYFWDo+BHaz2zGj0ZMLtIIrSJ6AbskkgjRqIbIGajo3dt9t9uz+CTi
UmwFKolzE9xEbobfyBIGfBni3Zx2gSHyIiVLhH2Y6jkfn1AkQD57f+Xy4wTeaYe0sdLiWqXSkGyL
YONQx5ZcgyryqcN9odE52RsFb2nMhj2VokRuxRNg6fq98wAEdI/v6kTNAAN+r7eYhvb9IkQVXrr6
ECdSlAVf31Dek5KE5ZOxmUlZh9f+zy9ZpFK9unJjLyvq4Hm17ri4RV+zXBe8AdDbeI1/+dsVUvS0
kXTFJ7V/XYNOpsNLND+T1/QcklujqRtC+FUA0FzdfiTOVGg2HT6sWZcp6Jpp+cEzDN5nVowmo1uM
uPu14aCJ7RpEEuPYRy1Dm1rBGPT+rvjQVM6sOhex3fjNqjuxVhkqmoz66Q0X/dvS7ymZD2AaJZiK
n5o+3ZRAjX4Sz9ydWJ/etHXliP1+mqYtBYqnHn34ai4kZonYj6szmovv5yvWnJxkKEhZc4UT7Rx/
oq5aJ54AolC1WptAda8WKeX82QODwh05BNGGdR5mu5DHV0u5A+dO45UBFLlcDKPaTG6AcayJuTgn
iyt3mYcqqgXxJPXQqPlCettBJMWcf5ztl5dSYdbmWJcyZfFmg9ClltSWnZ66q9Y93Iz1Wm+GMrZi
1IdQ2QXEHrep+XV+L1seZ+8sgOt7KUgqNaLpkumNP3DSVew9t/tee7TGeZsI1pIM51NOT7zAz4qS
EX9a6fu2h5BXazfNSPEcio9k3rHVxE8APLnAqEiAbHfS4/YjBw9VeCaPPSBaTolZYMisyP+MtNY0
QYZbUHtm6WoyDQRWdAtgyPWZtpo5ihKp0GnC5qKWYgztFRAG8/dbcA/Tgr6N/fuf3ShSizHprFs3
H+Ioa47AsPkejjX7EWwLDHBTaQNLUmbcedf7a5EaM4mrEGIn1FlZqD7BEfPCTaBu2CcBTr6N10J5
eTtFGlKzRj3F4Kv+eDwumF2LkxElBRXEgGZintU4+OT7vCY45H4f5MM1yUKyR8SBkyUY7d5VPeBy
9FCKwkU14TZ0hrLO6XrCcTqG99BNeX7/ffWUSlfDpXB3b6s4hcT9w38cR/jC77MQQpzoQz61cfZA
esvxZoQyi6luEYhUAUtnD+eOcTkGPfMjJSpzQs2rJaNAAQgnHEJbjJhYCjKWp2Gn7zO2QYWipUyp
qhxX8U79fBjVhExOkm59bCxSDrjXfBJyfZ64rSkXZX5hrcMk+b9xAgvyfwZuzMM3Z6Ti6t0pdOIT
TBJKjALIH4dBj4/MAHA0cyNWUled3L2Z63AHHSN5gJKuLvp0ffw0RdSjfw4Dso2MJwkR50tyEW9b
T0Bphktwj6XSZQ8my2eRoqelJfxsNNy95X2VNVeBbxoGMMEvQVr1ff3S4RhCQqxvsnIh7TLCFlm9
PM4LdUNcitqjsPEJsfhl83vHclZe+T2+nfn9r44k1MmO9QRp83nY+QeeydpKzrnweKKMN9XoVLlf
wR7ZNBpe0fiGoSnExf5xcRgMzutaQPp2GOPINtjTLUpgWN+uIrlE6OZ1gry53+LNialguuUZmmWU
46tFXBJDRbkudmOHGeUR4qbilB9/5yXYGFUAirQm8E7D7ovq0nyaEY/HEFzQxkGUmhVQah2yO57d
nxCxrpTyDf93YeL+ULJPo1+A1v5Q0raQhjtaDLKl6SfFI25+mm/CQ5GIe/xGMiuv4pSrCoTbnunw
eKAzO5YeGfQMcensjQzxj6GU95s18n9GQm28KyEaTXfhGj/Z56KlzUutYs43E80f3NK864D3rZ9W
OqWQLbNMVMGzMLwo9p4VFJtTuBRbBaE6A50es9YCea+XM8Dnd+bYm7a6YOTu36uyjUuILqK5x77W
FS4y2Ulc8Lg6BONV0sxBdCljGvS+ir+lYi5QT7t/6qoink+dlORnwkUZ0MW9Axxg0DCVUmhCEyw3
VxFgrXfjuEWVX2p5vUN6SymzfOlQANieL+NTmYi0M9a/30AcYX2uwZDQzvaI8Ny60/25VpgpiJHH
P2WYeHPuJ+eq4XXtIOHighlvf0vue6nVyJCSaEYBOV/IgM2kyroB/SvRBxC9Sx0oi8P/nLML7Hxk
GcD8LTAPV84Xfg006zkA9BRU7PL9OlKi1hVHuA87fOK6evAjsNqGLyQl8I+OXEgWAgHh8Ys9u9BB
wZzq85XBFE0L7D1bWd2nINeoAoeixHPOZuwqtvER8qzVvKmDctWMKQlaedAxYDecw+wLNNNmPkjH
ekCfCu/8wGkKSBAQZpmSw1XdF8MF3aBFrGk12qXEWhhj3I0cYn4A+UQtGsDuj2t9PIA1VRZV5IIe
fp5Bi0BZC5lSw2PTuVCzcotLmRruFHxobs+MjN5x4251XpFJ0oIszdicinRWlfsSzy8h+SapY+ST
cNquMgUx0pHUEFKDoZZFQAhgh6mSIsp6rkN/+NRhnDZiXtWK84YAiYvHeE52/4bsBvdnf+0HgHqv
6x4wgY3xUOSo/WBpakBt0B01A2bhjLjqBLUhW2cZOIdyXJ9bAE7KX+9snE8nVBsgYkPn+Ym6hosy
RkPeOZpquYFqwaAYstcNTZZD9oEePmcyyln6euiDlX0Lej9dafX3LWkcENcJaEvyI6jIZLAEsN9N
Pqfh+G6J5ZARU2t6ILuq6R/9nslkqvBWK2VVKUcizFGHwm4dor82YlUZVkmjY0hHKbmPWA5HsVoh
2oDldcWEZXuUhyUn2jERYy5tqig+wwet9YcAKVCCsul6KMFX8knFo3xnGkFPMWZ3GByCiabQmPaT
RXGV5Abm/UBfGKOZBl7GeHFHesFqRTpInnupJiUnIbdaCDVrJtPn/yaf5wUvO3+9EPBsJGiMUbOu
Q8sm0YKYeovQWEYy5a9XE/Ur8tPvw875Gr6qLAbGU9IgMBj9ioUgsIsKvH+0i/Zjt2igFBNf2fga
y67mIuTpIQkI82IHKTSD2Jk4canDHBeTIfvj1twwijCWILDKzH4NouAfWZCuSFmtRYrk2SeHWljy
DxqcL7TrPWtl2Pto3PRPe/od/7aRzRxRwwM8WdWcoD+NBireIrXSCoCFhrieh1wR24oG5rS/W2ne
20qwIx0Rtf3+J8leRkl8uaZeqSYA+X2lK+DS/Sth4zJvGWExvj6hawvXSRhco4UX8rL9EEP6V9/U
J3R2EEiAtfVBhzTCkukbrbKEu0mJVm+4CuZzHES41NVxRUU/nIgL4NYLOPCQ61m0ZFIC14nnzGTv
1fdn05rMTdoahdswx+SiEuPub6c+fo+euCOFzXj7C3O7xy9r9SkPaB73n18EPh5HMJsNiNMCJ0xc
ZRkBRoQdQWMfv9simTwb5ETrlrLIKOHlAH6CveBE8/YLrj28K1+hAVvByAlOSMxpyCp2jZDbuqjw
E1i34t6aVB9IejjMtdFtSmFzFn2Sosih2Zcu+DI6BoVwson0HMaEyZ6JHHB3tKt+i2xp37wdD/sO
6b2sYwW+7bawtRXzu9f5xOOzE4jIVvUnxx4iuyAhY79N1q9P1yGONs9pYuSLGohbfchWz3mktsmw
20I9KnlWK3l9SMkeiNusWQwBoniV0wZFh3trE9K2FmBOQfuyJ77Tuw28SVO67mHR27TtFdNWhwS4
zKPZhNX44B+jHHasnilUzrj7m+EssDtUdVXRhxf8Zuxi9MSL/CNwO6mbH5Alsp6bIm+gubPqdeBs
0Y733mQ3CB73dZYQgWLewPlfaXngqAQjBn4HtCKpfRVhFxcwdrnejXzc99yo4oNgqmkzbE89TcoN
VMabMgBylpNt8M07ycA1O+Mlg2KnZ/ORHjLON0pMjewa/RtUUdHZqREF4+eDlee5X5KXc0JNVoJx
T8XnuMDFUYR4FT+HKjokfn4Ybhw9r1n0hro2pWgCS60izwJvwc1m9SnRyxyL18CxkKUe6Q1qH4oa
R+xksOjh8kky7HVvW36ZpSn7HrHX3C1paLMvNXGWB4WDES9DrnVFdnPRIcqz/1q4ThzMgX6cZapT
XizalbndAT4pvHNN1e299dDQFH5/BM4hSyJifE9t3BvvDYncRKNN4BEkGIserNkO65dCFZmJ64zY
06JNAlJzzfeUWeTdZOzjSewkdK9UARcIIWGIMotCpUk21rB5q40TSkGobqoGDxifn6m0uj6NWs6l
ksZcOhL4tZuUowWgTxuMJg02WTZhmEaMmc45hTRaN2z63We7qn1LTo7mZSxZnlrXSIiyqAufufL4
0K7fo/LisRzn4ynYSalbyiontZ2pV2XWw+msCyoqdWR3mNQGDJS2DmY8BEgmHCONUy8mEEEppKl1
EU1KFCswntXRhZcoX9fXCONxSYSTVLOjNnpEXQc6WtkRzoWWW5hz0Y4/dCTmVeBqnR57Rr1WWWuO
hUyZTaPjllfX8Irjs0RYD9WIRWl4nq0F1fS2nvM6cE6u1mWw0Vl1bzEJ2yobjKlm0L2SuNq/R+iP
dPJlSo1k1oboggQ0VtzmjmxenR0KDxuLJcUqUqh/h+x+GhATdqZ8bXklzHEc7FsHAhC6zxPSnmaB
TWuE/fGPRx3pTIy7oEtX9vKlbd+B8BO6tVAmYhXEzFlETR0KiWgearpifvGi0wa7TiHj78Bh+XTZ
NCSTH8x1r4I5gI3hJOQhL2JSq1iIDSl5NWlSlJ4qiQIsbB4zZakvjEB8U2jwkMcmp0s3IWQtYCQY
BrI66UO2LBbebjUU63FUc/t9uTCogwcaqAIaz3PSLyqbeIzNsP5y6JKDhS5AlpqS+/SxQH1Fb+vG
lhioAgJMMD5MEHrO5f0VsOlIUNFgNeIhKdnlQ9LWS/T7kZnjJGX5VNJPSlJVliclYUlCi8XwhX36
Drb5cjna//84WDvbNB/wv+j0FX9PSqC5qGapyflYDQ2tvEv4Hj6UXjlxoQyseFXbBmZdZmglfIWQ
COWfXrLNWgEwfzXDge3Z0UzgjHlKkvqI5w+SMHu4nixbwWir16Q+vlV4VjDqs3dcyJmmW+n71UXU
tHAmuZbxBSD15csniFV0n1aldub9bvsL4zn+q8mX6xhup27uwKRrtJKRdZCCxJ4baQycyGbx0z9P
0mQyg+6hBl6z9awad/TICRZsJAmvlEHxuRi3Lzxhizo/LLZeFzs71VTE3ty1SW9Zu22G7z/Gtcd2
QzO90/wgi//p1nHFYlDps+8erj7+q0ScdbtC0091joEIhHYSsolxfXGcE6xfowPUALMMJaPmOZ5D
lzydRIDuk9e8CppxwnghqvsRvslWeh0nobFfEQqJE9UqcLuhC4T4Z1h6RsUV11Rss/ElRVsbOX5C
ED8lbnBlTb0Na3UOGc10iwOxckwZgLYqgfxccry3GIOBOISTTSm/nj7KgXhzmX8S9n+7EGN95N5b
wCkjRX69luuDcyQe4zM4805a+JanQ2QSwfWkaByIRjpjG0tBAdp4absC6iVDewQMMFsx2u0xF3Yh
svdLWThSLG0oQLDn3Ep3dOkFRBuCsA8jet8rWuGZ6xtBmw6Z4mbylQ4+nIetqjdgk3BL4wut8DYL
oujvKqjcQazwpUj7oxRYD2WaVjl6C3VPj3Pzbvho0A1jUi8OxBGbhNc5zsYXxGuvhDaWiBBWDvGw
BnRn6vXYhnN0CW+kDN1E2ubLDJK4o8ZA0q+CAca7MA2bTl5EXbgYYYeDLZFSaBmFfRVFUC4TiXno
6NzCo8p8mqTATYq0eUWo0AOvB1tPxBaEG8/vQy3WHQ9u8KcyKndgAyd1XptnZoTbBHXKRZq3/wlo
pEWj0xCc8jKtJp0vfBUnTXEfC7j8sXQ4A/ct/fJXGBsF0oH9IhEsvCzO0hNauI3jMrBQSYYjI9sg
FFK4EVswFxLuipyDfa7cohBkCwi7sQolYi+a4+sj+0zJ1g8VV96iGNHdxI5OAXW+xC+i0A3CAVH3
agt6QOadPKD8PcKT8aJD56uHuLmYUjWYv9qTc7jX84edokY4f2T20m/WT+3NWMwnyt+qnURht59Q
yGRaTWl2w2DYOK3SraVz7DAbMpwDBHECJe9Ykuy9pODc0mmHDaGGHZo3P/NSN6Ace5/2LRsq9qQ4
knT8PSeiWriwj025ChWCWBZBSVlquoAxKgS0XiSxMQrazChlco1RWb+6q3qQKwQuyByZ3jPeIksi
2XzYlcHkqErrSwbHTdQI5jH8UhAodm77XL1xWjqLpFn1kOzAzsVmD2oTvIxgnsnhCG2hRBuyW7k1
x61uYCyQQKoRHMLTDYQiF0sghN4OpncFKupN+RYFPGyTk0B2H/AqaAaPw3GB/tU50UX/ws2B4usu
MKUKfcEa0IHW/80ZWep2HoFnIoRIBzyj6AX8vWHuZKcitwAnu7UBmqEiTDWX9FLe/mNHdM1w2b3i
eZA2G4yREbtuAYSUeGWT664+12td7/TcW2aTnOvCqjGwB938Q3RBNd6MBI1X+E7adPhDuc2qdPqm
EXMGWKM1zP93DoZqfiYn+GEh4tPbEOFaRdegi/HwFDxPeKH1gRk5ihQ+JyOFVeonLyzamkLtGTzk
/rfnozuyPrG564GK6wVDUsRo5LnMCvsLLSXiMLbLTyi1QAo6cgmXn4Uzznc2glMjqn24XN1AoWA8
2ARMARpSQ0maboHT2RYC5c0kXhvOWXEfD0HOmtN5ZT+U7ywbJUP8NGPFtfxM043v+jNV6zIioszm
+arGBOVUGS/9vWpK+ZOAmZ4VfYhhqoRIveACDzlJvpgxMDmXwoh5Xh9KRnI40LL+K8YC61VDHkD+
UTZRFzVVSNNFgn/8TVBcqY40RrUlFDyyoTQeEt+7HNqvB3DQpLT9j65YfB3VYE7oXZ2pkAgIAhM/
gEEj+P62Pg3b4sD3xn2iGZBgKN3rrSINwJrp2dmcsOivU8bgEohi1fK34cigPmR9LwjjYaQjKyJB
koH6oaSsu3j0CTPc5fHnkip3Gfuw3IOwxwWwg9fYPG3hmszRKIorwYvRLqluV5EthEm6WeXUOXL4
vdKXlLp+qNlbzWP4vfty8JH419vwu05YwnvNQZ045TvKqUZiJBh4dpisZ+eUIgTvwT9NnSmupGrc
PGIzVyYdmOQzJGKoctY6W9kV7sOME9/O2iKduCInXKSW4+P9nJd42BuDnWhngyS+ugndCWQxneMS
o8IDjFpoxTQkpfJfmE/YVC6MoNjGZPmG7AM5q0b4830QkKr3dHuXWRtSTPhbjtr3esiuNTVpaWp1
WcR3RRe/5J0b/ZTn4MtbfqltkFK8/jNDXumv99sddv0cYilgXNDw4u6TMmhxaFYxR37fTas4icax
a4eomhNaEz/0nnxpSMs3XOlOvbwVMwwYSvhjScj/J3s7gIjJOXh/6f9JqERqN3mYvwM1PruWJW8f
kxjfIFWHtXoU0NlZm/wFppT3i3MlHJzLMriNh4BC2gaePHyPCof1PN99YMtbTEBRPFhMf9nBGkz4
tNlwj8nBOl1926YBFe3+vGqsWZ5aJJqX+VFiWtU9XVlZuZYpiJKx7p9wD2tM2yFizWSkPU90kIW5
kbMqo8jMWSLFlAHjqLKwMLX+oREok8S/558PxB2XxsZ5rRtut+M11FbUcXRYev4XQcE2gtjgjao1
bE2C0AM9nHjxyqxAWyR4RM6BkuCp6yEY0fL/galCztdTVMn8IYEQ9cjaXkEr8eWmDWy5ZT13CtM4
P6vLMhg4CtrIEk9IbJIEzLMZXAzC8ovmFPIWpoufKSFIccMSWeUkbdBtOpzJgz9CKkFyPIIUsOS2
pvkexgKosmLAZS5WBp4JU2rzvs8Je8LAQld45Z0aXQG7b72hYRKCOnP3Wn/hdbZqI+Ijxgg43beI
/2Nsffjkx86xA3NDd1zNWG7KR7SpCdU9U0g+IbB95oEhRtQA2zbOd436HLAuwMa9TiIn5fTY/kKg
mI6aGHDA1LBjtRh8P+a5DiVv7DERAeys94c+L+K11DJr2+/SUk6rBodOGembs/PzqQGamimZwJt6
3s7IDo9z7NngJAgU8+58rGhz6NfmycfOtMQ2BFg4lRhZ1BqND6nsVbA+iZtm8XT71PjhPzjfauxt
uYfsSS+o1TAGTNqv7T0RvxiP1znPi/6Lg/X0sLM3gVeaR6utXceftPvc1Ar6/kqCPNqUYXieZ/da
XowP1lFVy9CFC1HE4POF07ZGYR43n/ZxQjNRYmHRYveuds8flpuuhQVbnHg/cSTI39MxVVWzctgN
5SNm8V/R/a8UNeaJSjV6PnyMKUQg7zcUTWejm8nN0oTKFBgCEFhqXaQ7CyxBE5EQp+5oAGBV8BoD
U+nk+GSOSUi1x88mSoCCPTnrPGP4asPyQozzDVlBNmplQ8qiNSIeHp301nS1oR8mXdsGeiAoNP7I
1lQbLYKy3fEWW4L6Kr1cR3C73NzpQ73w8MtWB5UJFRnwZmwDPuJ9NSzOL0xa08/heH/ypg2tndRe
eaO44DVGkgL5gtw775KcfV8xI3qOis0kUgNu+ZW7AMiARxwTugQDt2tagCo58CaIGmDDP69Dgr3w
ddLkCorL0+a0JF3CB7uszS++bp6TwK0w9/FkE4/qviSNWqf+G+XVvbwYDXd5rQBeklWGz6wpOFvt
w+MUxgzgZmyNez18HzL9zS+TB7sRLB9c6zgiG4N00GU4T7AOHq5gOvt1CQRJIOEI4BHfJQVFWY+r
Pw2X1v7lVs4Udy8El4/SazJ1Jn/7/08Tz+xkEnUtOcuctIlBOGd0h12tN6HyVuxkrgH1tBzUAOGd
3GP2VJ3VlehszRqZM392+ob4oPCMDZWFDZBRKBOHDAk+99FkreLYLpsmuPyYv8ACjM3Ldii002q2
sXKzgu0QY/W/Q8hlIArij6SYGMYptqjkk/bKAzUKEFFSHQq0rypuUPeFKBIzVRt+1gcYSN5wffSv
TBKyuncWLJ/OYYmkTkO22FfFJ4B5QvWgZVgIqB19kgI5Pt+vAplvgrz7Ce0JUFyrYTqkAICRkZ0F
UEXhU006ZVCSfaIVcv9enrtn7Aelbv6Vmie4UbDvraVueYk66wrcOi4eeiTy44z2o7/84xIk6DwR
OOoJ98F1B70UzE/MoSZDK7j80qyyaXm9b4rtDQlqGj328iuw3dSase5XSMwNIoJaPuzeBkCDlwNV
Mgr0POKQBpG7kgE7NTCjggpY/XJdyaSwv1Bgnguhtw5BXqCvGuVnOSUA5ROPbGPl8wKs8CWaEZKt
c7hR9gB5R5eUXtvspjrbaIxMQWSZtyQ2/+Mi+JQqqBIb1HqfFL+Fz2/bELS+uYTKOKE3XtWepPWc
7Q010uU6tMSJgKph+RihxTehD09D20uwkzQ1JV9iy5eFJjGGH/0D/8vGkaDfv/OMfOYn/NwTf5GY
lmyVJSjk4L9brN0fqWcfcZNuBYXq8y2wtFn02JZeEBPGLYuI72TeTFQ/TnGuJqdPFC/f/P7fBTLm
oK3TaPSHdRbuPGVKCoQBoA97fUbYhXOzL+qAihKo+uxN+/9xhvbOsl2vFOTUnow05nxSrkJs/Y9Q
clDnNQpWL2Ltu5pyEmaVw5m0qGqCNfZRft/xdGP1wvNNsXeX163XeLdiP1W1OVRDnfscyNrmEcEn
DHuUVB9DVuyRCKbs8Q6hahM3zqchp1RvB2GK0gCcZWMKgdz67noW+o8vnqSzQumjuDl5Au8bkOpO
k/irXR/LoZOwjHjARYvO/45hbKtmnv5ieDkbqQ47WUqPXn0g/ynTdLKaH104xVXNI1ydGEimPt3E
u8Id5oWYWOiL5uL/adNRrxGnHtVhN7CmDG/APkm882nWNLMXZocFUaBWjuhV7WwRk/39vsSfInbw
/jVSUceO8Kkz1/XuCZPMD/vPwQ7BqQBUiOfqgaes7OMTTG4kPlKn2cHh5mko1K/obQOOJjoVRrWA
1LMvV4JWDyGx9qDGQEM03Kqqyk3jWtJdel4Hv1Gya6g6yzZdu/7fujmFvxIa6BJac7PA8gkBBxqI
HOx37ySw3Q7jrIh9EO7Ube7yA0Gs39+o6SQ89esPST7gPLtJOCygruBsy8t0HXY3XQczrSHoMVQn
hQO/a80m0ImMXx9gFZoIjJ6HjNuJY+L6xE78dOOMMsBayA/E11GNJ/6LaqYffyklQIIS19t3/pBM
v9je+FSLfRRMFKXoJ0lQGuVvdKNTEBbsvlaSk7P7AY3dYIGrob9EeMc8eWZam7838/eSN9YbUiIf
6xd4HzeSAxUcBJiJ0YlqzcPWQVXoZK7AWqJNvOLVNT2nNp1aHG6BHIcgDYYfNfDWaK/ANwo3JrU4
6NksCgIqh2WbISsRkaQTw6R4rgBIe7dQcGpKoczvM/5zkB5tFATouoFr7fLwmyPsQCBKOckfbqNK
wFMFQApSNYfFOOaJ5G9EPFNWm2xx8mY0PhXVR15M9xxBrkQKQ8vLzpsl7kXjnOM7hOmMV7URrWQb
cpLkl3WWhFkIx/aIWrJEuriBfG/vWIuoWHfGYaou+uf2epkkSEeb2kY2RiHlNDfHT/MpcyeMJxjF
1eOlHIbx2fnxtydeYmWbP/BHOQggFscUm8GYuSLgNWqkoXZ375shgt0kBMZrDZmeOAqRa9nwMoTv
vHHYvVsxXieTSgCgZ1LawSYpZQH3LocOikMGPowoKhqtD9NeEw2ehuiLLIlYf0B5P3xwtyuuL816
OQhLVFgS+nEM7rfs29AXApfNdx5VQYj7h2Qil0P0+sDlcwzhZYctUILDmHl5HtqIY97ixwMhJXUh
WCSC6EJ+fA9x42ouSh4WOe2L+e0wcnQRKwb2G6WmxANIvEbqFyxvmYxjY8GgoHigr7T46/JX1TP/
xPJ5ZR+AXBu0a3pvWN3kV0r2jNe2PFSqPjn/ZOwwKUosjCmIVxwkBgDX2oWShd1HWGwe6ZoyJELE
XJz59xvmBEH8qHPz2bV1NKglGTwO6ccrOuGr7r9B4EZcECrDNRgRq9R12tnNuI89m0U2JMdP+d86
r5w18h8fWnUDD4lPD/d+IW3dqx37513hiwdmieolMq7jmZSkytmowvwmeBydOQwjugXOodIVlZCN
ebXcS8H5bhHCyvgUFAOfWFROGA9b3ifURVxPU61mFO2cn/3xh+TVHnWyAgZMcTMjGeX/Gue+A8cX
LtgfquNeJ1geMXVLEAURNm1jtYkF5qWcrsFxxrAMOZkfK9JdCdkIpb0Wkfnn6t2rCF6WMcJJwH3c
9a9YgIfkot6lWuTXW9kXxwhUqCRkAd13dDDRrX1E+l3bAmRkcH1ta2A7JMgDqVrZfdH5xhAs95nI
uyhzD8uk1sbDBJBnG0MUWugoomTjE6luWjX/EgHA9BoYbfonFOecyOTF46fK99WK3cT0oIXHJwOp
hPZOGkEQioAXUZiHIcDZQVPnAmxgCh9ysxXK15n/wKyzXHWs1s6FXfawrRUP4PlQTm58JM8/8gRY
vs7mazLe5Ot9esgzyIuMBSu5uN/DdicprLYNKiM/9feS6Yy32KY2pBt9BkgSbzLzCOlMTD0Xj8aI
D6wt8lU83lf+gIxFZAlyz1PIUVXxDgYle+BohLVcaCBaP3xEUAm9a6f0frYYEqghIBe58fWl/wVB
HbK/hRsZ1nBKW87UTcQJJnVgG79mQIA6uMOhAv5GZKiSEtEFR1WyojJobpqeIhpZjrLEysXruxZG
BgkUqsOZb/D5CnfTybDnJhFO8QupX+jgzeOkd31VzX/TrvlX5f5Lnsbx2XJ+7eYM3ojDA7rpTvLl
v8nrMWcWEFEePAhr6kAYOFgtoAV6mFOPwqJGIKgFXvxRpZR1oUXI5R8lSECvyqietsAOWXCmj2T5
Oz8PQh6gMnIKiQutanBLj6Xi2+XWqdtidkRTW2vw9mE1K5EbEM0zHX6pdy47ENCRzCVFK9R9bbeK
n/WNEvnT/zCIUB3x1SuUcicdFM7n6alm4DKnOYd+LZjjVqmJQu7AOFfeaJs7nEutuFCQwfpvGIsY
uqwD70H5ZuCXLM6SuwVRtL+Y1T4YL9qAFfAASFP3j7oNZ+yczEcCz7vhDowsPMC+4ZD816ctrOmM
rIj3unNHpG4SG6iDvC9TL8ER1Tit6K5LL3yOzii8gn8PjXS4Y7eknGcOZB3JKyTtd9g+Pp3gBdik
uPZ9Ed+R7KiVfUD1nPBX9Ejy1n/skFe4out4x7gJP7ifPer8YTTlfAit1wj9eGaERNDEkZzkkPkE
PC4aoFmuMtoQvXrikXVdMNh+XPNXX5L1ZGDU+cxmk5+DzrJotHCSWM7evxEYSJxIQZzZgAed3oyO
dKfb6QlQfishaZzrO6a1T5kQcjJePjKDpYXLzOosV2QNC2aMBdb3TDyz7ZLy/NO2L/c46fBPrnRD
9v/TVqBZhkIvelV+sEPkcTMPB8G4pzkzFLDGYlu65v6gPtuLWaaNt5D8xBCw9p8NmglYXxS83hkn
ibBgl2wtSuJtP71beQfTh5AO3v1qAtgsSiKeoI5QltbMT7QBZgEElLE5u+wwWW5z93OkbH2kgbVP
jmc6j/tC/QQkF1lEGsJycAp0pwiVaHkJ62jjE5Nseqc3XCFugAT/EyTDgCSGLmNXD/iZZcF9Tymq
9eny87+HZjGxo/YFi10HpKCknMS5u5TcdVvz11y9KLN2iBQM7B+9CEafq1cH9UEYOtlFe+jXdVjC
JGxA3td14YkCssxA5uWLengVKoqQAyq/QxCM/26OSo1ZwkZL748HYu4MTxQTFgsX532btimT88Tp
p1JtAyQRdwJE6Kqi0SyaiacrwPsV1swbaTnxLKsys6EBt7ko+cB/nbmyZnifxoggDL8XbaFE+0Y1
4FwrF+51TFJZeDwec9AX1jpQgtFeCEo+EVVOA+9K9tOGrQOcfoYjP75BSUX3g9eQ8b/UR86cIBUO
+EQfSMfIhMBf3ZlfrLBM9qzfbyWFE9g5VVZAVqFTH0MTHIRfbPx7ORrMhUuRGqd20QOPMSdm513f
l/83ILkcUOZppP61ySn7HuhNqywa+rcY19sRwm464kzOJScx7uU0WkZtH4jqhSb51JkB8mf+wNOL
FxGU/6g5FV/yKDtDQIpAMfJ1ksmMmv6UP7zb30ovaJqq5WxiCfHNueBHRNLu8jLNGruPIKRp6VDH
w8Ylsm28e9sDms4ohTUTjTAW59o7J4S1NjcdCmwoMknRTHbQzEe/QEV0SUEDVWYkecYEHuYG5Poj
lCBb12D+u4E53q7JZUunXyygo/XKd18xKqKx3kctINnZ2+RuzPFzIvdpo5LZqZOyp5W4zFebwGKP
k+7qVQH/zWncK8ATIotxYE3YkSlnZ7lvYZWDmOngP0b1+/g/jLGWhBHJdVU6aolM9qyqAS7uDL4q
MzsbgKINcPDocXVAlhx3LgitlvEcZ+0p42LaiLFrarrk7tNqjT9JhryRusrXev3ZNXGayyRGOSG7
g8PGs/uzr+qrx2P0pP4Cvn9cLKj478tvNJk4Sl+HdP8+f/MabA2oNfBgPXvw5jg2D5QOQBo5i3hy
9kW6icMVN5GYgdk+0ANSTTweQYgxGNx11zoxVqqYB1zckfcN13iSR8tvj0moptjP8mQ1cTKELdv6
2MCFZi/Fv+Uf/E082bQ+exxRWezxpjDOqehG4U9ayOEQmsiR7FtukY+SpqW73mTNOfhgnQu3rJnO
/r6QurTjK/wSp/o976RC5FEOAFOGY6ZtWbtOpaFFlqOBIvN8HRYWMSkdIRSjFN7r/YDZeer3qSj0
VKmO+V/koGkdbfm9e/mUHWU8qpVERASN3O9wiTc9awNIHzItHZMRHh8VXu7rD0WZwBoasE5+I/cM
TAlvAdk+bVVT+8wGl41NMunbdbfvHUMB3EKPVh2iA2bVwO4j62hmJpLVLgs0IQ2ymqCqfFCnsumA
cZEtQxZHWFjVvwfkDYO2cFeOG6T/iak85ZBlbqEFplgv0MQRKrxclqQ/1mnPyfK7qI2Btr7j0Z0a
txleywVncsdnA641EeDB/I9sBZ5u2tWmOgOYzlhJHN0FvOF8wAOorLvrD2pmtLQEkx7YtuDfBwmo
gLsXHhtmlsQXxnkdhgZOAniolj0vud37Xm5JFBmz9p6t2zhUVyKmVU/lpwyTw34VNdieQOgisQUk
64jZk6Stkq5bIFn2hXtbIRdSmr/9aI8DG6yhSAg9qowKEpkxGT5eFeGipluTdL2unnldbVAkc+Gx
AqAiVNdlSA3r2FMzCclk/R1gdbfQERglUFhtFXnd0T/9LJrEJb/8RCs+Rdqc0Ojf559k5I/Dp3BY
qSAZJr/Ws4c6YZg9/hYS5fj/KS3ANx18hDq/0lJWvdGx2Sn8c6MGmKuzhALZxKqVd5JJvsCM81jL
4C4AFJyeFcArGEiOoMA4Pf7OS86Yl4A5GgdB/qn3836tHxqVvtzzlk+HWSVsC+spKjbLozlZxODF
GgrXGNNfSv+3McWLG3QWny+97UpKhtqo/QpgyVbRkazDnlAnEnBEJQ1Md/n06gk7pe+JGkN5Z5Ba
CIe8/vHfWnavXO5a5vQ57HpDW0ajNj4P/rWHMZDhPEqf+fXlvTIHI0YPSpftLU27RZFaFjqW/RRu
HiU647xcPndlFDLlhR03CMf3XnRWRzzgxBlLFcpKv2pFcw3mc7TnMej2k0ItsWLF+ZpPSh5uUOAp
pPKrykGcGEgQrZtQ6f++pDyVIFtUrGpGDvuAM0oUt4bgjuukTSmRIbmOD1uNBRCVR8bzj5FtoIeq
ebmA1KbPr+2K2XgmbMGYT/r3ha1jL1lN1eBLuNGP0fck9Gprb1hasR/YGvSl8rRWPJDHK9bYT0Tu
dAMboWpctIifc42+wS1+IDiD4c8Agf9s0jNOacOiAp2mmuaqlGwFTOJk2zdWSHD4PUKbyXSOlhaZ
3P1sqQYZAcjKH3iU4lY1lE8zy7H3EN/2DhCk4zaTvjJaAO/oo7D760HJMkZAWXzo0L7twvXZRa93
joQ0PbDla/OnsO/ZCKuYL9fI1cykTBZbDiowTlsARdjn8x5+VwiIYdZIykXS05myZBnhmKLTLVCd
DjraDcnLr0luJgC91h0GAkpET7bDfL6NH8lyGoeWull3sXOucMlb2Y9x+jU9JKuvdywUM5QXs5Pc
IlkaIQwYIK60wgPk+kdgf/QhBvEspMr90qegbz12J7wrDovmq+AVQEbOtpxREes4dDNDgdm4oUfS
E64iIoRrPpyDdsDoC/caE6ioyLeQaPrFBhDWxZlNS6IOvzrs3UraGNbZ5NUunEqPHDDecijb0L9+
mYZ7nFOKuwsdiUslEFaVaytmibmnLD5GKxiIzFYI1WTWXzNFZthFTHZlLwYBIRDNakO/Q8rdGJng
r9OE+r50DxM8E/c3mE0bDJD087ir4vEmiJhVJkGJAljkyy3H85rhyXBkhYDJFV4niEk27P4VRJkv
4aHqX3mlpT4AXHpJxQzN2v7JThoiHmUkyVk5IdGKRwmRNAjjB9R+AzTKtBgH0MyBOATP7FtX04B7
cop0Z/wePrdrQUVtQTzGNnbxg1etAVXivtiJhFIWvUR4EnmexCO8jLN6CZa0AbfMMNLDRSGsH/b0
gWFjxTOv5cWItDwD88qNH4D0n4zAe2JG1yVf3enVHdsXmSBf5HAFmW+P/QYmteOPPXC/la2azrqN
t9MAVz3tH/6hioXPfVERoHmgXsXkAQNqNUwjF4jXWBgDpIgpKkCLJK7S579p2okRnbKUe4dnCwEM
+RNrDRO8CoIkzTgRSGBime1P+qajWPz8UyEJNVzWwvWojLkCYpNZYsC1hKcmRsMRoxAPhh2zGrLK
ddC2gR3mhHGRzDgTze465C/zflDdX/LzEMwCTLcPToqBCzmwP1s58i/+nehX5lnVXd49ujX9tlLn
orEo3A+yJDoZNkxbSawLTYs9b8LoKSMlondohqU0MD0/zXMlmjHmtaQ0iMoEE3YX/SNjtnrPiX/m
VcWywNhnA85q2DO1frDYTJU9pX8J4gR9PcSe6DLTrsIvV1uza2xf0iekGhkdV/n5pinNI9geRAVY
3PZeD305VBn0wvmrq1Z36UubUrMbJiUAGazf1CJjrdBJAuQdckSWau/cAZd+b9s0gYObur2210tL
eM6hAQjvY7N1ZR0Y/leeGChXlcM0/7fimtwJw9zIbMh/TFfFJ+vf5FvX41MFv+/r6OU1pL4/KnKF
6iDLWP5TcMIrmL4vB4muqjPsxU6GvvG/8n3ibVVaBNIwRkNUOShQoBmPaPNZ+5B2E/z5yAmcfYgS
VJvxzSFjCg4wi/Y7+ySdgqFF4WOycIzLRx96rdPDD9x5+ujzvujIynvHHngK4LZk+WjBn9Avf7eb
gTthq7rLFvE0XK0TSBq49DLB0/IEbDNFU0YiUTFmfHGLr+QdREeHsXVwjd33gFpnvjs/Giv2VEjU
q8ilJyIsgtwrOo6OcfWqJ+OUgtD52Hqh0CnYdxv39bkknwjvmIbiQF9rmJrcQBSTZzePIMFvpj0P
4cXIHvCGFKluCwN8rGDNXs929prabraMFJ/rvjmb/BIo8C8lJDMoPv7kmsft1+fTylhuFOOQjGcX
lU5YIupyqxYih3Sy2ezengn6gDP7shn/TBqB7ZPkz15t0Hqz/Ozo7n7FJAuk+lQixP1JIA5XhteF
cX3ruNGJeQLVVwX7lh9DFR0M4suTlHzd32r/xj/NZZ3UQ5ZfvtXL0HwgrqhBuLE+5Y+ac9bkyJVX
rTmfNL/aTP0CjIDOWhZEfVDIreFdyQ5W5RdQoBIRpBvRHxHueIS/pJ6QmQtS1R/XuMp2gLxkoUaA
sIPBXSwcn9EvE5uIYlYEqkmPA/GpL+saDfB+v98o1fv5cLeFF9YXD8LC7rjNsPeJ2z9d267KmeQF
zhfuEmU2moEFft1K6gkWc959HJpHJu325cfKChg0eEhclmlUS9l9ysVPpbHS8uAwLOfN9yfdjw/u
0bIAMe7TJ+IaPiWWW5GT+crDLriJQ2aOOg5Rjm1vYJyLfYN3zkf3+BS55JjyPhKHEbBWo2vP/muy
5YS+MUvyQrxE3OaetgOXbpSSIuCf2IkHYAS0SVWDIl2u8P5cpJCtORAYjZGIBUDdOdPx7qqj8Gby
KOncbg7YLFLB7T+PYgOq463mQw+iLDOS81ze5DBH/4gS0lt868dZH35mYntuj70rgjfC1ztAx0L9
Yc/9r7kEhxKRDhnLHhrsc1HYJH8DNdSaaGsd0hfj6vmWDMwSzTwTl9DgQmemIrkPL6RxG2lMEJ2x
Eno32ux7hNE2OV0hDmvj5LBeuCOBM2NQy+p9Fs+zqY0B6vfdCFF98Hq/algs0mTXyflB+r73gdxE
xPNxOqrqv6Z3TMwbzG/C7gXRTHxgApSDQzYqltaRbXUwXiLP+86/ovbjvDlv5PaM0XT6zl6aHS8P
OpLGIxUnLURtZ6HpMm3GkLamCq+GHFxUxNsRij3Yyzyi5Ef6EdgOxbrYg6v5rDc2F395dgppogFj
x6MVstYVy6dwEk6mM4Eo65J2FyX9n2LMNwoViml2acX5YRovaZukkGMn9DrEe+XDDq1Lh7pe9eDD
dnDWG3z71GDJ5qt3ovsJR7l2UWlQcvWBw8fvIKwghOB7ZdubDlJEbXsSIRRAkBY0II9vn0Vxgtpk
F1YOqJ3MWnglzHBoSSUS9OOEDu+fRYinQY1w2pGFOkudSZF8rk13RU1Q+CDhVQrXQBWABGRPS1OS
e3qdN8I80pcfpv5Aqih8BUjtVx4Cep+xPy7veF4AyF5Q5xmfZdCQy9b1YsdD2E2/A6Uvx+A+Gj6b
IDDDqGuOwq1JWhhbDGuBgkBOFpuO3aZIj/QOZryVHotaeKRPO4KrNoZlkubRqxQwHN8JhI/Pmnn3
HW/EDVO+UdQL7cOfCbS6aKqzjSO2dXSzRSsCp2DlKW2ZUrLONw4JfrEqruQk2uCjPL2QCktTZtNj
ouccaxiIqRxKSVJGk9xEYCXhGMMb/Ak6V/tHQkeJX1vtx7F/kmDVIJfkkQFfxzBMJ+zbp4sR1/tw
PkVZ+V2DdVNxo1LmAIhZ4o24MD8lvQ7TIk/YsED1q8Z0ZBOpQj4in8ZT+tIOhSuBf6iUSpYoMOqk
5AQZM5RlFd0e/q9UP4Z7jyF8x6w+jv8QVVpk+8XRWyZKroWMpqD5YMbJUAn9NIHFqcMlDXzaaUNs
jtbWHIqddQZxrKaF549tqe4FFd6H5musuOoD9J77zCvhMZOkKHORI3Tek9cr1d08b1R0v1LXiRwO
XFMJHuZBSs7aDEvMldIB474BPnXDr9KTDfBZM9ZFUNV1xr+Ic6JJMg+UAnaX67EQxpVAaP+gP0W4
52d8yzI3E+7ZD2AcFjLaK15SCBIMoDHxgP994ctIdPm6x+LpChHy1f9hsAS7W3CRmjDjhhIoLb4+
dx95YzRzFxn08xQPXxcMxLFBvKXt6y2Q/ldS7BsDI/S3HoWWA+hvGf5UeK6S+cBqkuyUF293kdUc
hiU1lBZha5VqOJPxvGYjr+dCFlJjU4fW2EnMCzzKP6cOMaB7A45dcYZjmcH+9ptDU6IKIa/Pbe8A
zZNvQBTU3sgACPNlS+DyryILHAY7UIr4lq20dwxpj1obWnZZuFvScpuENMIs7kSPY+OHDV/CM+wl
kyC+y9o9GJpl6AgWVGyWJW6boMUzAwkcowR+SzP2TacEYEMfeOeB+qcJTCuHM/M+RQ0Evptwyi/K
dOQYKeuqDd8V8yo9LehJmjfVhCHG43D0zWKEuWEI7OIFn3coVMdj2gnfGjTxsDpybdkdsUrYbsiL
rHi/NnbF5f0t9pXm//Vm7qs/g7R3a6EQ/x+ISFHg7ym0JklM6Hni9YfoG64OOZA4l3Z+LScYrxVk
JDDMYLXEYMcYTYrbwSHk5IallGWsmBY35bmvOXL7kRfUIAVTkF47QThiE/f0iYgOcJdUP4AB9Mau
JOTeL2i5BakJoNOA/yAu5eJ9LxUmEASmo/2jsS/BG2f+ZboWZiCEYg17z3Odlm+lf4FCaAa7fUIq
D0boqUSGkdfsBlBLV0GQNzjrBPBjqCgj7lQN1Y+x9wXQALkYCMC3C90uPtdI9QCVma5oAcvoZQc3
LIHgSSk0YcNcIsaj3lg8qClvfUZm3QLA6OA0dTpceBhCrlf4ybAc61prp07zXbmfyncF5j48fVa4
qv9zERGXpByo8hNLOUTY8fe4diHLY4d1SypuryAlyVv75pNw5H7/FpTwqob+Q/NnUTL+ntu0QWzJ
52SV5mEt6WqY+5JbPveXYpRcJ6RCCwTDuPAXLZGM8dovV35jSbMsPGdDA3B/HmXiWcKML7cPW56A
vzdS8xLFr8TWBKBTEO92GW+ohC2qWYfqTiZUp0IC4s12IlVbD8Qb4JCX+lY53Lf57XVR3rEhzpNP
l0WDnLn2k0fKywFFohpfroxP9jNusnn5pG3Jjxk5GxNIDvga7Vas7aBWlk00xb2/g2gCBSnnZWnC
Hc9D3X/qpIFmFa7XOyrBbx1LL09u+jv2zmLRm//xXp4v6bpDgnFqdsabsZwbYdKbOqPxd8gEfy0J
Vn/qzVIny5wpleLBT3/sW7e3qdTpj0NyRWO2Xzf9Zbyk+vipBH5G/+u1U0zf6JQI7V4S9F9vXgS5
iC0w1HT+AkY204VW2Xw22+WEVhzFDY6MB6qypjfaVKCOW8qnkv3Rs51DcKujgvvwhHRH/el3coOR
9xRwaiXc5HU56UmgXIp062m4GXdSFKb73apTZc1uMYuNnQMmfHJhak6efN3UPyQFViqfdgoHeA5V
/91mjYfqSUz39g4J8q75AY9JlPDo5+nB0a3Z+aeExA6TnGjh7msHh9O6yTt4uJ5De0HS2wFg7QFc
vyLPF+MpAB3flfViUe3yNh7iEsrdIx2t6/sR0rW2D49ZgOXq7hWsOblKYgIOTep9UBye6I2lmJIU
2POKwTzKjR0zzXoCxhNzyl+CHRm3USZr2A58k1UDHDNIOTpYpJSlSearFG9lZ2jFC4B+rL2fb0f+
ggTTMQ7haILvDPucNTifnC5TQMUt215f/5QcxLRzwLRI9AeLrVGtQCjS3/wm4hRMWEn1zerM1tlD
Ay0YwkmVpArsOaMxTwjW0xH54xhPPvXkEnRQ2ZQ2tnLiRDyrs2teCCRLnMGyMvCA9FHJQMMSSv9s
bBnS2ZrUZoGVoPOmnV2JwGPuR5hSQDsJ2/UQsZgdYhh9IIbVS7yjzHUQ+E4Eq0/71ueBtXNlpFva
UBMjCj/FzieCf/UZlcPzRnK473P69D+Ua9onzsRl6sM2/fJvuHxLyeRPeHZ/7uSMjpmYYLcGroWX
Cp/ljisps3N3a5/4blA8gbvkHc/CzN1xsf9npUvqHQMk2ZXWrbnX1wA3R3TbmgCcaeA9yuOdOrFK
6gkZZ+7qcmRsD9QUCxkxTp9BtfGr3lpim3BmpTvn00OjIn/Jc+gzaoFIz6QQe9a1vU/pgRKy7kQW
StiYc/cHKhsyyvv+Qev54b6uCSbWtcjO2a5YAalxFVYB7tedEwrH0pek09upd5XIy+rD6cwmWKsg
RPpf5DvaB45lGS4AQnO0E2Pj/pQERTq2uJfXZypIAhLkhklleY6piaYAip4tmLy2tWimVKi6ql6x
HLkiAQhY3q32wTDo26xarf8m3T+PBSUcvKYT2ffTPlNtXyU8oBM/X2bUFCZSpZgs7Sc7xuz2lCTs
97TCx6fqR9bVddHghF//10CKnRpOTYgzXwLH/cC+wLj6tCdH6LLNMpdGadd/jOk2OyUmLC/Qf0am
5RRCIjHk3J3bVsRUN29BPJZei06wCC6f1jAIkebVOxwVnJeF9IRTHexBxye/ZT0sRX6dr3tOWxjl
qrSHoJCMPUk5jwardkQZICY4twT6L3PmiSySKfLTfMizR/3nnhcrHcY27+9zkALKBWWfU9BURMgL
QfIv3R8WGb9CnxaHK58jkEJoCeven5yG+ojYSBkt7rDjzlKY46fft9b/im0Zx5teWSN/hj5bEeUB
CZuYF97WDnQdk+Y1YhU3WkgEoMqrTf3PWO5IZFQCf4flZBnKtTG19SaxVwl+6WeXtxyRkvSGaeXL
ZurT6E/mOXfX6kpvqAi1/ZtcuAQBu4CStjFTed1oJqa0cj3QHEa0YM6gToahAG02Z61uG5CgW27g
lz4OlGs/vSgF6WbboeIcON1MIXtL1QiEBOT+8A5rf6xvZQT/PcPBvAJmze1QblwugmRUcYKQrkvN
ws2XIPsomT3TfyPD8SAMf7HRqrRHOzhigOm/MDyUqn9l83BCkGJLCJmxbYsFIKPc1VPpj5gyBeeG
d5ZgxalNk8tuPdtfj3FjLAg3t6lfU8tFimFBigfhzrvntEp2SQqXVugFEgJVDLrapK3ZcXFWunfk
Q+bxycsGWgi8vtxoUZhL/fAvxFvRZexwCJZvd2d9GResWl+wAAQJfAmK1X+2dSWzBbg7D3yvyH+O
0fqr8tPselrAN2GHWj1G+eS6x2tw8ApOeqgp8sUALDK8NfFLkmJFT3zbFBmbVMi8Of7xu0ktgXTt
K66h8wS8nlBVhCEslnCL7RaYxQ2kB92JlcQqrILu0UtGO91cmze+Y5YMYouXmNdNOjN1Z1PsJkay
3ZJt67UnrKnxeXGovP7ET2EWroW6Gx4NtKMBe5r82oC3CQSZOfhO9MXI90XhhVBijY55m/HQgSep
CoBWNFuLPAJe9NLdjRiIDsBwgAnIhftNE+KCdnGpAYU3AuJrA9MkkJHDKdqXf9SdqWbypUXpRIhw
wecx+47rEdnKEwWWT78KN/pp1mFu0KM0ug+e5ZWLjy2836IAlkLJ9C/CBg1xg2wg6Zn0K92OE3IX
ggCrm1VUFPJwHHbkRQDIIOAEuwu0EPbXLFe6HFzGFnAY3GEwisu6NJpwXXnxrZWjr1A0XtShdTFh
lEIPUcWAn9ThL9xmVc+48EuS7IuVTgc0DnfQZHLnVkWd7S/E+ZGzgHkW0UvL2s2iz4xl98vlgqr1
21/jg9U5lSm1TpmLy9H1VBhizwxj8DywABpYZs/3v2x2rUwavAYrqcOa/EOJ04dKYgNbgI0nJF3D
SNR+mRrHTHlCwcU0wkJi7dp0fHeGy9ujDV8YaJ06QzGzrqdGbnQ4rMPystd2eCLCxpt7nRkutv2S
/dY+QcMnaPxdMxT/BaXwQ7kFGBpJcMUFqn2415zRC7jVxpsIaNdnQw4zO62wSXTJlRF6T+7uUEsY
wqgKlV2rFvhOcq7NXiooiI+z5y4irH0zkuvDR0qXX72G9i8j+LizAUIQnz8W2to/wZo/QMOSnRlq
SmH4iRJZt27a2SQO3xxd6x9uOGO1Xml998Y1XUWqclEyT42+gqVvd/ST1pmlAF13fVDvjh5lE3VK
0sH072ezo3GtU27QzPyWpLfTHAYp291ZdLKSRZglrAYpD23YgY/NmmREexxWOXdogfuOkcgRCuJf
C8WVHRvyAZn9zHZcfvc7inzB79cwIBEwyyavakXXv6Wm5PLsNNXTgnEydunQFIzYJnwsWK5orWLL
Z0GiuEP3z949JqmTJwC2UpCLNNBLzCprWkHvx1rXiNBFP7igvnO6nO3q3RldCj3sI+pXJ/m4QHJ6
7eZxsYsOJoS9/LkZkvDOYDM/DVYhDHTIEgaPBflY69DJkDWYvTM69JeGjWaX2ZQu3W05lA2iHGI2
2XkqJUX/37cdx88IfqaxisJ28OZT/ItkONXRT920lDsoqElBJ4kdxM8+WLFZIC9wdBW17MAJHsgV
WOh+4d6XybhCefmihUBsaNd1klEtyXaQhBD7nB2gLpDhS4aGafkl1AssdKYf8IGWaEOLpHi2HtOm
c4tf4F6Hd6QDU7bqnyF+llGHDkCSJI9XeVLOSBRP7mRPlCGJMLnPkl8mrmCDukCQRcav7C5ylUQ7
l1IfBlgNDpm6yoGGR1cO3r5zknl6T7TDjdBQjZKwvagrqZePhHYSv7P/mfN+1dAQii9lxNK4X+aS
5ID1o/I9wSqCy8j90SkIxaUhFVpYit3dDv+vU4xTSEfBaRFLl523dnqsb2E7u/g4pa4GccH4bLDO
S4YuCRL+KjnlQ5UxVHmZuv1fU0gaLMUbH8s8qCzFNQcpIAtm0r13LQu9tpw924faEBsyEsamgpSq
P2SCwbuEJYeJjdVYucObBd+z4/3t1AuF9lxkAp02APjmL2slsDwWooJWFqZ7G9ZKV3gJY2NxUJxU
MYHhtWzJQvZUzTIMXQ49axN2Et840HU/ccb+QoPyrBMv3jjWmiVSK9uqgRBZWzQ2jOkZANzh1p3B
G98r8NR9qVCWGsLypiLhZeVmQvx8TVSh70TeuFNuWTqQ2AFV3DWBxZBXXInIqr2TkNr8QTH9jrH/
EP4iIiUnL/wOtNriAq+hFJoP/rINsaRwDIfiHF/usugM+pcRHuhZjsvZKjTV5766s1upveEoV3AZ
S5lwNQs0fek6uzjaCc09gj0AB6f4rKs1mZOZfCX0jSJ4bNdx9CCEYEAAa54978On+ZozPaW+KtJQ
XWTONpDm4IZzfKic18GG+uB5hYxMPgx2gdLntz8tAthUc3SIsruLpGwKhNhD/51MWTH98R5Dj+zd
nj4Jbo4jKksP1jSYNpxBD4Bf37UETrgBD7edD1yz4jXFLiQ0FiCI6sS16fejq19sy2EOcvLJ5PiM
HYFniPNDkS3KAH3K9CoQarQoW2IQ1E4b0zi9Pqnmh/70195iH5OJftvzPVHkfTLVPzpUl4sq08ym
1J2WN1vtRnqV25Pyvm5k/BJjLvKP+nTEEgd8/BihJMRNUt/RPyOV8uyLiDVHddQ6b1yvNtw5dUUG
vugBfYLCG9Ix5Cc7BZuYRQCOQML7dU+WSjACMEVoIGmje3HW509ek6MXB3O6hypSwN72aU7SQoD4
Jg77h/AoiwLY9T20El6gqH9XAGzAYpdSnXrpSsF8qQ3cWSNQ4I7fAd5Vz2vBNJd4SYLKpqeSB7Ps
yBsMWBW9XOaUaf9NtnM2P+kjdKlpn/TDI6AVelvEe6dt7Gj35dxEHMYiMpksMF+gFzxP/ouky/XI
0Q+zUqzphXCgG/3VygXmFeEfkt7mOjs95ZdQJPt4YF5WAI6xM8r/psafnT1trjfcp2nqVbiu3imC
XyyJ6REghPcocxOoRhdRYEwpFCwylSuTdfCT6qc1QlQEX63fcLzHGmDwzeMm9G++tUf556r7yAFP
3YT9D58SVydrk1zpOpdjbowy2riuepNmO7CHl4dChtv3utbu4+1RNTgpHPiKPPSH4uVHp991ZN+7
xFWYy/yP+l+tqZ67TP2haFuxQ0QRc2viJsJOK1Wf0mP50satXmJDzRu/TZ8kpq4aF7sV4/gcZWx1
X/P4+Ot9QBRJF8cI/bAuMeY8yuiobkfkt+Lhjwk86Kz3/kNNg60LPnTnXUsakOZbTLww9P00iosh
6V/sI4DG7zcak7Oc3vWWZWvcIxX0MdjLMC4L02YDMvXkbA8xBTT9sYYTbQ0JwFwTmcDPxVJpvVi9
Z4U96qUp0OKF5ZugzXTE538hBSTPBseqp7omuiRB2keIS2H99O80vtlHpt0TWrEwcFyOgSNcvGqy
FevcsKTwSK82UT0kJfQRyQsiH2gLZCUlUPUehFfhS0PVS8A2D/2GxU6xumtqO3rAentw5MyZfVku
MPUcCEvgxkIEEq2qvyLFwysCce0c6ymMYNdIyp7Xt4900p6SdEIe3HYqmIoVDS6kmTi+X4243pqS
JG90JzgaRO7k+/KMZRn4NLAcYf7+XLWxhI0xQb5cJOwa4hokS1EtN5zvgH8Ka0D28TM2TtEX8usA
jjTiSzcfCqpwmU5HY9BifFR3t7b6d75Z7QMnFdZxcqffzOyZXQlbypALrQmpoVbii8OCQR0R5P09
Iu8YxJRYl7TIqLM6+AubZnXQN+UyCJAwQ+ZfJemVp5dgzi/XUQYxx1FRJxilF6e/65rO8pKAjTEG
ZEwE84SonT3dJqqcSue48ECLS8lkRVgXZcjHcxzfWiEF/8frSqGg2o6garSOwxY/Fwe74ftGeNud
ttRJfAwLIS8Ygapj557fTdVfjoNgSc4QnBar9GDNcmAdSGkPkO+M2medX4fYpI2yRYDwZrest+P+
XpgRuDCvqPRqXYoSS/Rs0QFoB9MUp24XptKYoethpGdvddnAgEFUgn74awAh5k7F/f1zXqHqev9E
EY/yqolZiykGOWU3U48NX1wLm4oTLLvp6gV/xgKGu3ZZWsWIClV0ewbMjw84jPzQJrl24cSfJN9R
URhSBAmjWQCauWk3ZS8s38U7MivSaySeC+CixbPl/GTQOJzdhHRXGdNB7JWzt2Y+xi//4oE8/3k3
SX2oUXREBY3TZXI/7jypAb+TmvfcWU76fy/RmxKmzhJ9fCL1MUIxgj0itpO2C8ua+p91roHGhXEA
WS4COahdqV9tLLt3SToy0bYYmvFtglfAQsQ+JkzOzls/3DXJ4NTKmsLGOQe+6JpmKAlXEWaatGvf
7mK6oZ+lJANS6ETd1J/2hSJAXluyQlUwCWfu85nAJ1q3XDpjT23p3Yt37/0GzceDTr8Zfz0OnQcp
iCVSc4CTTmC89878TWzJG5psVtIQYn2ZBxwKdF5lDanuAg8wJOTIkhUqagHju8RkwkQAouqzONzp
5C4I5PvGJShvym0PnEKBKSf4xg0nHAZViVqyHRguOF0gjAxBXSQ+bse9koQmpnGfewEbbp+h+3jY
9JSkWpjJw+S0IOOwzcah2/2cGy9APrLrvckY+qBMX6sabJLtRridvTQapnCyVpiEXtj6ydQEad5y
5gxPo8fgO90DO4qkWKuAV+/kmMlsnG5mK6CR1gXBQJujwh2Dp7HaggZW6wczOG/sybu8O6NDiIw8
JHQVSTjZdkMTyRv66vox4RT1tnv1xsvt2uQZK5XSaF2OOXkV2jVlFFxqEUhBTKyaqf3VNhjChWcZ
sMRv23IZX/NfajCR3C+Ozck50S1W1EWkMPUGvCrMPyqS1VbzEM0PRt1FvczRBOO4PJ+8P694yhx7
jkW+3/6uGPIOPRdTvkaJMeuSNpPv9nBMi0nWEiPxj96Boi4YK8h6SvNqABAH0esIAVrq/d5obO6q
6TQ340TXOWnsHX6VxQ/OaKc8A8yBeQ/nQ3RtrWkcckfU9bWcRTokykrukIS/Wqy49BukEndXdlqS
1bnyKc4B7k8uTuLGzC9WGpX8CHsfB7mIpFPJMGzO5B1fYY8wv+gFrS0APWvD77IulRJ1umOLsGY2
3KXAZxsuz0stv1+LI6I3YaQBs5tf0HzumMLfRC2mViqMq7eL2fQeNRcuuh4mYxgw2CguiDcF06F2
pcpmfDJ3jGxCuU2st4sU7RSLE3hu/kjZHprPdUwDSqEXK+7qyiopQ2Er5eAonkHnMEUReQYPLEt+
mm6cXebbyfG10UZps5d59giKE1fnQNDkCjXMtiqPnmEMncQMWJSd5fyXopSIUNCw/p3jXWrb6dlT
yJ6w8qfGVqdXOeJ+DYpWrehz4yOJ4+/MSKpSQUPWu9O7cyobSf22Tn9Rs8SBbH9cIVkqZf9GzWbk
N1jt612fsVWWjtJlaRhMZwV0lYGcgz6GIBxMtn2lc5pf/+u4vrx0dtTEwHrvRZvJUZt/MAv3CkfR
TwNnb/frpFM/2JMvxVJ9WUU+5DAbY3+Y5W5y0/kMGge4da+u+kNlJA92Dt5MHETS1ichI4AaKLzV
dzry60/yCs5LAlIQMie2625KuJm8mZr6sceFsj21GsYA7KdhUJ5wR2O3j6MeZK9UIgkGTAAAIjw2
vrcTO9ECcwFkD7xJf7kql1oA5BMFznKUCiKpFjI3xO3E7WHuwAKS6xNjwA0p6KRjXlC30idjIP2V
wjXFjNwEoX3o2J/H/8NcDWBSfx1rBA5i4o0EftCea1Y0icHZvldlTcLNWbvIqi04TRkDAkxg3dnd
0+5nlZj/eI7YvfRL9+L/WK0dKOsnxW9gJYJbsW2zYLaOjn/LaDgvc6YR+QaPi7tQCN1RhowD6gfb
d1CsOmMJjFIlnggxNrka4GCEca2VrSCBUAHheCjp6Fdmmbt6kE6BXNr5Ns0bfTzE6hX0OCEN3lnG
MfLRyTjKc2y2qqLeHQBlofWXboumyABCsRyKD41dYttcYr7GdWcKncVzXH8kyH0VmvoKYWgBNE7e
Rh1j+rJvHJhB/dOqWuqFyeeyR//dfK3tRPhS1Nk3/zFCAVJv1jRDwCt0MHR1cbuRgdl+APOS9oR3
ua9+m82AZ0oBtydJzd1MuZ7BFtfDi4axMvW6350/QquAoOFkzmIPDwRDTGGGTeZwMs0hlnp9RlLW
3Y7ZfcvzpvS6DpAEu3egsydRcKIbmmShvzzYT/FbAZjcbluuI6xBC9np+uAJiCq7nWzpS0q8U4tB
ArN5BmDVgWIWRuUYiqxWgYTk0IgstqVhBl4EE9UJxLHtzupcAU2Rxt9yP0SAjPvJkzhD2kZ4jv48
OQ8bJCALwV5HFQnCYUWTY71sblF28Kpvc5bx5DOI/RCgC5uTb9KzoGpJklNdtNXXQT9JQPzaRxg7
LNQnchV1piqgjwj8TXXbqZymkWpa8Cfwl+uekoXOYwkvd0knN4hCFxpnIqXKbxUCAFhfvZu1w6Wv
FCBHvOboWkGNCOcaGwYUm5jBZ9XhV+SMArysVLJhJND79DaSct//JYvi4Svv9WH+KpKrfOreUIdv
9CYHJN4/2HWmNjCBDbs2oEBMxLDh5JUryIHCCpqN8YM3SVDPTY/lsSkrWT9ZyxrtRx491U9IXtHD
htIvfH6MapLBPG8EaSHjywdJA42xBoy1gRxTG4Jh3SinY6p46wWd6+EC2b+EKQl/yjOPcQA7wIDm
e5GPbYZQsiA5gpjOxEXOV/rpHI4z+8tQughdu6TWF/Fy4e6iY1vX89zdPMp0ffm5srYviTDLj47x
HPx2hAdVM2h6dByPtlf8Vxu8uE7NLwbxx9blUSJ+3hzOqiu4sLqG+DfxO0Rj2BctFdEJgMzBxgc5
M7ZzKy3rI/YM3kvDjl6KUMHL4HsvW6Ub7Rv3F6avDpIiawAjhVPttd9ZWrBFrgGsO6npzAQ6Xhyw
IT+pVDJPhrIk6v/0uEi4bzqSfQuY9xezP8E4V3G2uHCeYCr8AjT4IwM1OpZGFtn7y7B6eo9kD+60
0N8yt6tL5Yox+D9yqrnu/XH41ExN8jKvTc8oHGzW7OgOL9ishBkC49uxVd4yJpqUwrIx6HkhXch8
eB+oH/SLhUEnuc4yZautaaotortkBVzirr8iXuyOTbEWZmg9PndW26MKzpgHLGntZ82zmkiQPrHJ
4mnuK/ibK+0iYdKxDWxTfvPgy3fruJoaINDWakl07I3SdKIvM6XFnHTZ5d3/zHyGYpceOKigkx81
XQVCKYhJbfxl3aVtGQdqEH0IuqBt6TB/WD7tQJ+W3tXR40+aM0bTPuFYbgVZUi4VEDmFZ6V8JgdJ
SKl6kDXDV/xGehENK560oElqxdTtPoCTihj4yQrU2B69pbKj4T2vBZq4wluiWDEYaDvI6b1sMqJ5
gg7Cj/WY1jGifEnucDp5dow5fQGvM3G2IFIcu9zys9m1Mjr9tnzBQNB6AMbNjQK0Ty14Ka7idxiX
kevDVI7EceaVgO57XusH+k0I4/q4Y24LtV5oKqdXDaU9NR4OptxTroKIttTtLNnoHArjeaFWKCkh
GR7+wA62Pwk/NxTf8HrERkA7woN/KiwTpIjDjd9Tpdhf+PnpXP+OOMhudng1TV6XgRLdRq2F2SdJ
QamIiliS3ZTxCdO+NQJ5GsaJ7QPFPrMbmkGk7PJsujKabb5pit0xECMhZU2+Bh61U7OqCbpn4WUs
JtnWbdgFuvGuxZgmYVelIwEx1/27hAFcpV3nUM85yW0b7T8Rf4iiKbWdAAoQ/SU0mDh/GwOKdLBJ
LxwIn9YqIQmg0hLPUT3jafETYmsYGjR8HEETY1f4Puplu/CmS1BW5hlZFDE5tVaQVc8TgXEWv/WQ
RCqeR0l9MpCnRqPgDE9lUaBNJJLBzxUOceUFm/EeGzYfaweikoFBUOlujsSmWUaxGcZyxzHZR1lw
peNC5DvEC0kUgxhubsS6axMhXBpdnUlOtFT1Rf/JHaKJ6eYTHkGEt0qgeDIeDgCsbhyGSTTnKlLN
ZlKomy2egy1vOKZQ2QAFmhdtbafD2m7zH0u9TJZkFnnOPackp+mTaF8bcidkPLe2LlmhINi8ZYkc
kpPWJGK6026OX+xM/zU8vd8GWLvUmfri/tWKUb6cKfPx/XRredi+PsWoxIfJblo2dh6HCv92CTK9
UBS01pa6m7LrgLoACkNSYYT7p/DUZ6Ns4f3rvQ/x/wNs53eLV21OJpA20d8kBxj+LAyS+nsqf+DQ
oQT7ulTa1Kong86ylweECorZdK17+4cZW4vgIOhgLJpuusZnGyaVKvX7gJvul4DzPo/5MNKaW4we
Bel4j0YjsvsQVa/AMTNL+pa8JNHbguzwx7v2Gg3tolD3vvLf6oqYvPB7DRNmz1ynAjJ4QbrowvBZ
hROROVjl+/TztsEDT6lg3GpxETCdjOIZed25WXcU8QeLBMvYy8b2GMmDSEyBDEz4EGib7DbgLGk0
qSYr3Ye3iz1SJshTbxZV5zSMh7+WoQMrahLyS/C+Y80FTZ9xEW0lIsGpOdLFLojcnUAYQUl+C+N9
yyDL6tlkhQuS6BtyEzVAvemVpEhh21V7kxm8G4JrwlKTGJKTs76FnjkUfolH/H4PYi4JEUnFRU6e
ZwStytBZycfUonS6X0IENwGfnW/BBTNqTYgIpRkh3x13c9UjIk2BWrVTDkYAg6NL4FxRotgCOM2+
k/djnPJaBW2zbncH6TUozET9K9OtHFpl5NI9JJ3nICZJH6VAc619ZBBDffUV5sNVRp3r6yFewflt
VF1ZnvcQqIWehyYQEqVBQIPYkyOm9W8Q98vdcgT59GFHxMZWCK9rSZcx588pd9mQ/+hEngkP6V8/
Q9C4St5p+jDRFCNxDE6H0e0slZaHoniCNCTZNcxr9f1ifsDIO7yk90r5/XnLGWtvdHbcNykb+p9E
7nqetPeccwSmzk5fY2qHmsMvJnU+vJJP3oeArxqUZ1nIfvvKilFxP5Xq5WkOFyw7KLFcRqBfIkko
5PZdsTtAHl0GQKUiXwBvF+vEJ7y/1DHQBKy/7FQ73W0f3F3uBzE4JuN+jl61lq3kLmZEIuyYjz8s
u55jApq3tiyvhM4HbBOT19ZV373xKvsPNKGMY4CwQU2Lc5AblRJ89U5qMXhYEzW3fN0kWGFWIUNs
HvcvL38pOt0/Q+w/kq/NKhLmfeRP+QHqSl4ZaU1DrinsKU/tdupofk/CxCG8t1XVcoUCPY+10e/V
v888m/5600zVw7eYofoLi5YauJ6QwPOrqPN9/gl1XHC0OEJO4OHW4T/CVl6qZYGU1A/OIASU7v7l
JuH2l7svwM0gaidODHTSDoY7yYuQDhsxKUoOkeCQPoxWCIGVJ7xKxTP8G1RjjJXf79Seu+7gkDkx
7lONHwO5457tmDiEPeehX+V1V5omRx/N7XBIfSJGlOifaqmv/z6Sg2FFZasU4EnbYbkF5g1rKjDZ
JqE99MR4R/wDaORZh75A2u0zLStOoIEdc5av3ZPg6+1mWypifUyAeIdtw63Y18BcsZRvXHjhxAD7
PHgT0zBIXnEdyOMi+w18qjnDzbf8lsmRcs0Oh1HhRQUTfGMNxsx9wBMaSkaytI3gME9H/oZkp4UQ
R+tfmAlkZuOSu4dRTGsrERugtIEJZOZyzxuo75z+sfMS1MV7MEgRWaEOBEXzD7X9Ybb198khSngt
nqr6TfvMZy2QLctkLxgaNqIBUFbXBrGYR14mLqAZ7VavlkCI30rY7tmX9GTzaayFtlPs2JzivkNd
/Cch3l1uY3SUzu35KWY4+14fl6zTEVx/aFAE19rMALfstk12NYMvt8OIo1xUgzHQeLvRPXHdDFSN
dQWKSybYNRiXS1toBuZnN/axX0NK/pXr5dJXLZKOTPiemsfim3rIQpscxqJWr8ZExHleNlnS34R3
JbGzCSZ71ZmBMI8GStN3iueMcDnBdL6Mupyf9oBTnJYrPyJM9+HtGsxcVeomLSzRUaI63QFducrt
+rw/OEkI4HcNi4fcXugQZuL6S/9t+9MUZ6s9tigtOrX1pSYUdv72IwxS+mxC6ow/feP2K3EbrneV
b/AwFzF0/7Cx8hbh4HNjvvdcxNaDznjjmg4O0Or9kHKrjHodgaULMO2SRc7LbSsUbxFdEy8lKaXH
feqPBiNDzm2o5uMqn6LRLLWkNJlCbx5BD/Y817od620Pq6pczrttSoTOwx5iZelC9XJ7LQZaX5Xy
Y3Y1miK53C6fsvTWWBr06jjsV6vdLGJWtL8u5zi6PPCkJQvklCgs5ZdhrbcdttlrRRZg/yh7QfYi
hQgpgB+cQk+pHefxPlDkBnEDK8TnXdGfy9oys0MSi8yeD41NxqTx9fFkzt8QGcgYBCjrviLqxvRF
GjSWA5ibb8IrHi50YIiPhMpBbfn1sbf0DaNAlDXET75PypM/Q22gN6go9bxbxm8gaKTXg9eWOoou
rBvtEZRnqBZ2RSeH7NcUbB56WPzDf12+Cs8LqfKNZuKyqeyJ8We3qxVy7QfVNpalsFiDeeez9T4Q
Mn1pJ5yr5rNdr4fytlS1Q2sVLMU8Tb5Md7AHXQ/c1cAItWmgJVb901mTVGPgIQs/3i/nryH3/XkL
bVLedOuNXwEhm+d9DZhEt8qM0LbXXdgwhmg5CYnwXEbnwwtD7pYxW/fGDhEULR1UcfeMhQ6ob34R
5SYvjSMGg9vMAWSukXkIcdtgWVgO3x7PBtFjfNdNL1i2Btfs7d3Gn/BhYYRs4wdbKgsghgpF+WrU
+wDJhw+Sg5fe9jjkivG5Hy3Lcmfd8yBTG4wgYJYNlkv7RMw9vCfnW812FioDJrFCDsDYpkC4JTqL
GMuyy/Ku4sGNQakCYQVsHpuqk8jowM/5n1AqV8qBm/zb2/LmokkuM/LtQ/HqpQ24akrQ8+GP1X+4
BE0QrpXXptXc1bGBLBkY2MZ+AvyBqQKBWqbAz60H3NCklemLeR1hzCqueIRXM2BmDEWVx4sCNNDx
DUm6wm8gwWZSXxyRcf2zeML+8OqTwke09WDt7ufBm9ZEv0QermRVolNi1bgmO5AjUSOmT/+6QjzO
2Zc16Tevvn1GrEz5V2cx/P+xjN1mNm5eXR6RYqs9H8QegNB1bQddDzntqTdEaj2DkLQm6uE4YCQF
U+Z0JI6zSkSPCh7L3VQMDh4P19jkJYBTE0wt/Ks2ZLlJWgMAJ3ff9dubpn3KsCUJVrmMpiax5sFn
wX5qwVvTyMK+2yMj0v00FlSI3VJ/dY1KUKWf39F7QQJFDmAh2PbuA/kHWuQFfaHd/7uifPQTN34s
/4l6K1/+X/jIJ3aNeAknFap601kGNKqEjjoLY5NRFNdtWr3xgbtXsy5P+ePVUOONpx9gZGxLRQIl
IylzUXuavz+B5yqGQtk18mGdxb+TejfFjhvnqI182Gkw7fidkZZXpWIIlRoS3Qh9Wh4cZcZhrt7g
AIYpfEpnMDbP95bXcCj3sHvD6Ahv2Un7t3fDDpKQvTO3I3at4F+yGB05rscH5X9HyF/zheY83I4+
XJCzKd0S32z3CpU+XSThQVBOL8SUjug3g1JpagitO9nJgRmusYSLh9z38cPr6W6LatBK5WLmH97I
QXdpgiMqZylc+ggVFR+jBo4+yST4gpMXI3IqPz2iCosoc+YWFvB8lMY4vlMej8bX6oLrvqhRvHhH
XYyaF96Fo/aLiu6B+3s9C9IZYq3491eRZyy70/ncioDlHYcE0MbnzT4r9e2qvJaN4O1Bz/aB1w39
KjuePCeiqLn+v9kHR5q28susjVHvCc1MCW74nLtyfa9m9LoOYTDNnPDKjjaG/UuCnFbSxgDLJn26
wrVDrJ79MMOSGucsotXw0iKnrJd/9g5SkpU+RJJFX+q3kDKcYjeBvzNU/I0dRHTYKHW3WO/L+Snp
I/ybaDuEVJAbZZlAHE6O57kBzh+1ou0fSbtniczNAGBS+iwhjVh02JqPd5/TVnlIbt/SlBHz0myP
yI2r6xTfCCxtFlMowhiK+RS89thOpudX/L3fSmp+2hdn8EK73Ar4ARxuqBgzk3suPGfsmlmaD7LR
O/eBrYSoq/hcK819RsSAAhGgL6Gf32pBpoyCX/N/+qXXrFqGX/5vmlTJBah2mQpRqaXFMNqPpm+t
W/ZFZ4w+dQqHkm/49vRqrLTlWfG9LRA/hc5gQRZZZpAl0ssXOfBKUCyUMzFIuDjSx4VZf01CfHhN
ZUKFZVL6aginoH0VPXFqOWfE3Mf3I98QQhZTCK/lEbDOuJV5zpQbd6d2kdy2sRbLl4ioGzfO+QIl
AO7VNAM3rEUZcDjJv0QX9Fa0FL5XbpTIwAwGr9/HKuY1jD8MQAgzXPIexjJtXnnPYHuHXOU00rlD
6K9Yioz5CHqcta8NuLYpVBZxvFAKEfTkNGrC8N+gY+sTPktvUTnvAYTAayySyUT74hlOkSAeje9g
vRD7JMbUfKr7zvyUkHysfO1d9S3M8AccG+CjnSb8KM1N801exlU61q8/psouA9/WiMo1viWW6pix
AV77mTYbBk12d44iDL1R1y7UmAl7qqsHpAorj3HwtXrIJWxaov17+f9Fq9N62RK0JGMbkVhxKoex
T0s/XYjyoqpJnD1OTZD0BlPl/5knwGdn/qdGJkT+VDu1NUxMbyJ5+ROFqesj9IJpJHe9VITFpxa5
V4DgBtXIC/GDuPlZEZHgosfCjEJkT8arfi88SF8zwCciRUbc+0hrDkf6EYN8BdgC59TS1g/oOYjz
l3hijFnD+Ou9UzkqIAEBYDFI/w2hOzzWQ7yBJKdgdiiXDIVx0Q6yLajc7JqGpai3bggV9sK77EYS
rTNffg86BKHXhCdWOzPQeUSC6RwaXiW4+s01VABVM3V5PgXw5mSSAzkrOZVQbYoYzwkqPmMP6dfS
ZQVLfgW6Qg+Tsdqqz8iGNEF9eRZbVko9aprldKZtij9zMTN7QW0JXyRnKPYHSdTxM22c1D0WipEG
dUi9+u8PQq3sbQe4UVlSW5we1YXMlruCCtsn1iN8IQ3Lnvx2So+6Jf0x2RfNiADldwpEnOa6Syuq
GJVp/HRqtvLtxGGM1GkxFy+eg/2ZS5ssyMrjSLeV1iuWzAyJp0OEgCh1gVL9oQjESZwaNZDFxXTc
TNaOQIPwfz29Af1ywFIDPg9CK3n7li5njwnpwbyEPrveI0lV2E+XweHGM4533CNdgAYQdcB410eo
3g/11xts+a3zZHvvxa7MxiHEVUw3KVZmHz8Cbxzbs85VE2qjN9D1/KaZjdBAO2RcxW1DqKFzRtpM
3pltdQvbqqL2xiRbv0RW3SI6DpCwaT+vuOTx4QSDhf80F2DZP68pMS29yzhRXCxHvUZXHlC8aX1X
YsbkkyGY7pYsJqALEnx8YGs2Ha070bffjl/wYWJyBCqm3csb+Dif8Y2Jv/PWjsQ2U4TCt5vV3fVl
4U76/WoEiqw4Gpy2skgzFfDJJqcJihDWiPoDvPbNJACcTrSPusg+iNLJqI181JJs9pOxk8PmIl+0
tFYIdYz8cNXawwuJb1cw1CUNck1dgSoyMZ7dlBAmsKotwk5oCl5VVYKKOTsD28+snhEB0/yXL6vu
YUPTcinJPHl84kwwU5OSwG4innJpVcspj33yvDKy7lZXAZwPnKr1uKwZUWzlL2aJldPgUtbB8x0X
hnWbfC1HaJEbEJar9g8gJgfbUdrWEsrLV4RsEhQms/RZKzOemkj+mB5GXb6PtOJz4Jw11q5vjPT5
mkoL7PU6Xq93RXIe7ruYg5KnQjtb5fLicefXejeSfNniIUUcMccbD2kmNGvYO0MZNhQvvoh7LIW2
gWwikhqhtlh//7Mbz/Y6HiKWzZs116LO0XP3RHdhDMtFYl71saKVOQThmpCH+yCBztVLyZN2sWLp
eZ7dTKa6rJIlSuq2mPVQVklNdwHdZYO0w0EllJvcUsWKj93QXDZdSXG4xNCMD/Nz0pguZfpIIGbT
yIVqtcppYXuiZbA4CpsRexNIfpntlGQf9n6psXTQTIsp7DItcA/W4WoCi7E/MW5rXI4vidk7eKmB
VhUgcVhOzA9FmYggWiD/vTeziX38C4VIqfSagIL0AAGBaUT1xk0oddDA0S5C8cc+4bykzGpH82n3
ZNSn2ySKyxhy4Kgpwr02C7uHQUkxhEXD0R2cI4RjmHkflOnpY0sgYwNpc5SeLjsCU7y5eLJts3ny
NgPFTd1oRmrTJMxmDirnLidr2DhooitYmRaOJvKSrJl3KgH95rtAjDpqFFFV2Jmp7OmskNEJuXPr
4Gz7j799dozTiR0oTznii2uFVrYm02jD2d3g21Z1mtuKH42gyYC9tEiLK67DWQLMHCCw0YHq+o5y
YJSBK59cm9Fe2g0/fDTpA5C5vgfa3eQcSZ8BsexSD3lCBQjtw9gYxBDmlVbFPwREImeM+eHD6BK7
5zmkO+viWAVldU8mkTa7bnWkUkVCnclO/vZDDSjsjWYRI2EYAmbTURRECrktOgWFVltJY8Lv4Dou
8dGmAYRan1NvCrqaUp3SvttOR655gUrvSQ4BMuzhuQPdZACjaDQkpRwxQq/w8AxMQq38Sa05dbbv
kQm6dbSJ8KClHSV9TI9pBHxL5qrGS8QOjHeK0PfSCb+zdhD+GB8V1s6xSQ6I2vWaxY9BXawBJkgZ
BdJrKxidoMSNQ7p8Hyu1zvl3UWldLUJPNjk5yJebXPQ7xoLZrSab0q0d/6+AY1wHxoI0EFAd9cot
x25/nHrwQE0K2WSxDYiq2rRwhKR/RaTp69QjEXFoYIcsvxap3se7WAmkaIof2O+K+nLQRnXvF0Ti
Lp3vIjJyd+ME1101ENZvdlAkyHO3rFaX6Q6zNIFSXXRmcOtkOH02aJxR8xZJQeS0og+GZ1PMa/EM
7QemyNuvo76Loye404ynLunZrMnimtr0BH2PcndxAaUlZ6xeSU86/0S0ShAaeThBMblnDNH2ydaw
wIhQH23ec0CiqqJ0tLWK62Hf7CxtGbgBqcq16+s+nIHQhUWGAX2QtAOdNx46fH4dhPDSH9s7ATMq
1KHECUWISyVViNytC/pH8xIJxQQgOOLIVInWDe0nlfC1oKWEa9XzsMvDD1egsjlT0IaHqv8ULlOD
BzzhDHAbuh67qmD5p0hksfXXBeFfwLoifef1JAM3wrkvaFY/h4FQOwZhWG2xVVgl3rzwf9Zw7V6C
5u0Igg+UVWHzZL1LzfvF5aopBXDi8yn+1P4YUcFpvBt/61q9m7P09pJHSZQspavlr6b+IIStBXsv
RE67/MiswQ0atwn0yIOZ6KKG7JNcJhtE7P1kiJzUS3cLA0Um5IEW5ijQBUMXKtW3toScnHvaWxUP
Q2+CVsrYBErdHoZhe4iykeYVHosQu4ZVGjlCKJF32tLHmvvblJ8O0yDu6ei2qAGgC4ol3DrEzZcn
gcQmnaCzOBsayGse76BaTTRqnXDzOKMA0YSR4Q3X/e90Hd7S73LRZrEclYHk78urcXqtv6h8n4lO
AXMi7ESn+V/ElP2AfY50kmsrELwEAERPKfs9H+yeaZcxqaEOc9ya6+9xrCMCeGPOGgcuSbJ56zU7
ISmpvJDCUtykB8RxcoLcdVNKwXvxTamto3/y+yBCFoEx4ddrgcWntjDR/fETL/vs4nLZsaiRcjR0
0kjWxVypgLvzLArAlcGee3nx7229pVh2mX7bbbwp7zuf+O/zVrch2+m3+b5qdNM6V91+g7OlyAoB
C7C9TijwIKStDxIAw1OKxcMccJN5y3j7vsaWRb/kTnhYdMsBgby4oadBfd9k3oxJMlOZGWOBoiiD
AOal7dSGTQ77YF4jA5OCZy91lWmjKs8l6UzDfRR87CtBbzd7iB/DLXO0x/2PtaJv9MGIW0dqmQ9V
WdnNvYk+SPyUEYEhirk3j1O9Vi/tNfptlPRGO76rJcPtaDufg2rfRqZzjlMpADYIZf2Qj1z0jiiJ
3YaN1CWjIHijbQP0XeKBaE3DpE2blHYlNi/nVqptPB62B4wENhxbYSmYVyJ49n1jjUZ8NaFx9cXu
OQanR7f41VocbDD3Iph5PXLD4zkP52sPf9Pm/DG/34udwzMf/rzUpDKCUXOZD8i7CFSWna2zthkV
xS7tQ2WqU+d9Ui3ZLYIXt+rAkU+YoNPHZCV6PYsa4FR59kx9S6C+9r4uguUrFJtAXQ6eK0Rttt72
oa21fE3QVXnP+pr1nzaqvUV1vxXj0xyUj1qt4lJhri1xHnbfxgmOoTij1C/BScttf3yp38ET+3g+
m3bOvi5x22rTG6cDdf4EXVfq3mmOEbd7lKnuSi6b/vByNJhvui3RfA5tUt917Raowq/6J9REErS+
iD0mwEE8Pwjb/TTBawrjeZ2qJzEAI1CSKzAOFtx5iLfMvHzTrJt4g/+zlFjBUrndSs5E5qtuAtkL
7aWziv0vwOwX4PeG9GdGi/K05q99AKhuys8lze0qmB+0mtYj5Dnf3IY2dOrva94SLZBK3j5Vwi09
UiucodJBk5nPPEzLvuMak2Oj8u2LifylFqzlIEWh+Z6m9Ocx8fIHZG8phJ8NDDunkXmyG3xU9eNt
k9+dh9PzLe3lfNgiei2SnpORq0uIA2I/z83R8/Db0f3DVCYiIT9a6WaH0ZiGF+t2tsru4nNK8IGp
AlFOV8R2YTQ9hz7ydmtA7qN6tswtuteGaPHRERxGkVYXA4CYqSi6u1A263V94O8/VKJKGth590S/
WIzNrauE13ZPmi38HAJjDBWMUvfdCx8Ki0uxnG3W4YscwfmaumUwLb82OuxZDGWykFxnW1JfWfPJ
D4BwHBRNLvtBRttDMzn4leZdg+DdkpUQCXQPOwoWturdltoQicYVfQPtwCcEPTsaqokX+Fpr4MJm
ASgu6W1UUG7ckCfCNcYRNKgK6UkeMQsNEYRN4CAP5svR9kwtNtUcHz4SlegXWUeMw0/9htoEi1bL
GbAa2uksDD8Sa2zbb1be87UGV9T3LTF6mkqxapsbRFlx/QB1ea8LWK7qfRQf4YaH7p/t50BNFbG/
RL+fNsHslInQxxopm03KYzlHc3OhrqUPYHTPNwzj2dVQs7HwvVarsMgQTeGzfyGP6X5/IL8c8Wry
93an3aSei5norUfeEAH/DhY2nStE6593Be3PFo3jin2KhsADqd3US4XAYS66loQ2+9GELL4U1TJa
lsNiLRwUHf9XDirwQi+fzJHmD6fNejZZXNW+vVeUAnQJHqMgDOWVPyUk37YzMlbYB98bcWm4on99
VX4oaKlLBvexjMO7xBq6rWcgHT1JHatFxRGnLVPaA3Z8QUnqsu25ASqyXYKYPEjSFPTVY0WmZVwf
SG8nJl5IzoMUsoZNRhz7p/LDyAddU1Q6Zcyr/GNvSnUytHBlF0OpuZP8rrHZjy0s86rgpCMycLqZ
bAhy47znIQcEZBObGD5iS28iRgrWdiSc9Hthf1jnEVFIAJVsGcnsaVFUALlOSq/ZvPWQEf9KoHQb
Ko7UpyiHKGDVXNd/riAu1MiuboIInEdLtM3BAdiZwKFknq/TGtPsoY7EJf1+SRqXxEDSvQCUS1OL
jt8rtt74P4wt7gTtX2JXGzzHJ5tLldHsczi+YGW4RNDQAA4SAtIWJUCV1ZkHV0szTzab92PJ1KQG
OU9iG6Nyac7dGnNi/Cq0cyoON5E7/6fF0iPcmYeHcTtoOzEZVPqp8Z0CZVWLOkSy4kTFXx04rdSU
S7DlsUZbVOuBI0YQqQGbHxHY1d+FiOmiZ6af+FL2pRkgHrRO30tUhn4YH3BL/dCDL+/vGXXK0W87
Bb9BuB45CcsHlZVH3mTIbOIbDQQtwc3j94AXYjoLOYpsTI1+cTQZXLyAkQLNzDgKK5OHxHuJEnjd
6Oy2tO0BsYZfjS3ySJWdi48/024Q2bg6ETLfg1e2/vuRgZjk5Th9auoWSLx1yWlIUU2X3VrxV9Yu
nyG7JrJeT0QFxu69zGYMGF6LNjtxHc9LsCytaToAxIUnpZSaWDYVXIXucoySE8pgIc7R4LStpGjm
gJ/ZrA08/oIVqccjPgbyr82EmZpOZjpjr8pA/JvzgcysYv+msaZH9ePIaLq6Y3zVfHu59gBgZ/OP
rTIslaHgsN3VTlcUq0oUDKjDqQVlNVcSwlRiTmWB546HTKPLXzaax5ZkqXh65oMSEhAjNda2Jl0X
gWTgeIMZT8P9VRTKLUTx3NYGJgYX7VFfz2/mzc4P5h/ueaaXVrb7xDzK6fpZ6CytP9bwpIGUNIAO
q+1ULZtDsRXW+q6m4DDFZVZYJkx7Uu0+J40ySwy/XWi8PW5+FgvUuizCHCIb69xx858ZJBcY70MM
bpVpmcqTpvkpMczmhVhN/eaegx4gjSfeVvqTjy1mfSC1OFejXYWEF+sdHu41vhJFRwDeJh41U+J7
g+cKkwejfN9fS+Hp5mshDf4qchsM0ZEBe7E9kihgVkisuJytDLD4ByTgpal8k+li1MEV7P/181zq
cBLvQFd1BI43yV1DoWm41ew2TLuJC79WnZx49YJt8jdpi/wd05Nnw9Xm7LHjDAVVJLO+Wlp7h7OR
u0KawoyACovsQTpPAJ1OYVMPtGUbhC6svYVtvW55FeFEYvKnVdmOQ4ITV66hwgYAQusd4OZGNeVp
/UiL83SZ7XRz5hK0OCnWPgpPFDpsXdRB58+uR0ri7xFp/6jil+EgVXGFqq8OtQ4xvUIZ+Res0Ru8
RMrKJ4Y+J1Ec7uxMDVfrmnSXY/XOxmR6vSe+VYGvjYDP+qSJeJaR0Wpp7Lvk7z/meH/1GKMX1Q6q
VacHctthv0/AIjUx0VDpCgcz5Jxz1EQV/4X80VVqJ1eeBvh+tVwVaT5X92BdSPiVHQMX1YGVtYQf
zp8bvxWOdaCiwi+oolYg4wMcIL1C+Ws/UukMoEkiKVy/aAjRtGu3sHei4NfrwdLhfMDR16fyoFcW
SlNEZNNwrQg1Kiv9RUzNFx+ZsTc0449zBTZ/Heyg8za2PwcZ16ZdYjKygJHLrfAmI8lw+8J8+CaN
nGEvVAjI4kXuyeq5ssCgCI0TRhPSwwDBrg786/Wq46Y2rJyFuPHhVwTn57HyKQrWFnx0cpbvQJKx
7pONCD8oCdcO4R0kThwlCOH2SwAf323Bn0LOvlRBRri3oWJeyIj0EzbM/q4gfbc9dbiSvOIIK9Cc
jOcxzuzEWQwS/CdDhQtfWVQTTNF4n3M5dCByP/1iXtXJ8CaK0EgQfV7hsaxFqm4f6iKHH2ecZ/Mi
hCR5Yxdal2fs+tAEL2aRJ6EfNVAQRhEDXbZ0C0yM5Rg5RFWyYVq1BmCO5qJfFxziZ5YyYtUutlFN
S/1XABFx8VjCbh0pmAfRPaHXrafVBVLQJjnQwdciIG0DT49MIHu1R0CbGtoRR1G+xGkV7Pad4kAq
/QW0+zr7uB9CVu1cEAhM3EFd/y8uQtGNfE9DgaMKcmmx+W4+Zn+b9RlpOxpyoKQhqUgdaOdT7+zT
Im0NXaDxS33QJwCZGzrM77nLkFjs8VxD9Q3HPL2af24Rc//3JH05jaaYYMnoZx00SEjkpmoaXOu7
+TtFXIVBF605/BgrqGhi3eeoiK+1v99wjGfQMNaryhhlhczf31YU4ldigj1mwpf5kbKvHlBGKDLQ
PI5xT8s3Z9zLK6aD/ff52OkLHpq0scH4UKLA85rFxz++/8SWPhD4gkFDrjq/fL2yElHXTT83wP0G
oYgoH6oRS4guAXD0y2reEn/aHTN3jX28donY2ubjnIRll71S4KsSCBHXkGhzxM0ldMgIqZRPY3zi
DjqYqcdb/V26AGNqy5nwNFmb5JvKWLgXXQqc+yW0ZOIJzj3a4lkzJgVyV+hTTSMVaREP7l8ykfYn
GFoFnqIMgq50s/6KZuRno4oLLRPnp3wNMXNvpbyCdFCEUNC54I10chECkI8od3DNRMyq60UD/OaR
LKUrnpUatJIma/HoGBBJRbWQj+bpujOe85jVuxvW2At+nVu+x/dFEIuLGHTiiKiHZPhSrcrmpRkH
JK92V3311clrRh4WULO99UZFuYt45v3Ul3ByYkq3pE7TOynZkTKT0X5zs/aPR7SA7qG8T9fso7Jx
NNMriYHF9aoNRlgxVKLQcnoyGPwKtQizBMr/NdzGMb6OXnU2VAtBuqFcfe5pExqISG+H8bM0D5uo
MW2rEwgfxE8cfMrs0mKNXxSNir+o2oOi7BMUNkTcQ/AFyxShx23QyJubxz8NpzTIS6RH5eWwaiP0
LXn8MMy4CfdDyGfNeZbCCS16vUhq4eO+x2vEMaaymmQMtZXlkxwN2mNoE0GITrm3x2s7T04ffCZp
a4THyU3Zt2lIj/EUz+frZ9fXotXli9M1lG6hvRa11mKh1SfkQXqZ/Q6O1NywWU2OlNmsJOxOvH60
VJRL/pIQCM56cdc6AO0LeaxqmLWAym5xbKCs1bBLfkfBB6XiwxRFjJjfV/hDRwO+jgv86frHjZ9o
9cfpmd6Dc/qAMF1gaPEaHtRWFog9Q90f02Ka3uPnUp04UlsXRBPGqqxvITA2Ptnfn87f9yJ2uJpX
kSd9zqXUFKQknTJPZLEu9tPDwyMNbHXLsoKEYqtMxLmsjANOfrdC+cn3pUNqRR9+mVOZxEmZ1dlU
kImx1uCqKNy+CEGsSoEcO39iAljsF1/ywG88Z5NBQK+BzCkaDN6czatXO1LV2RXvpxjOCukWjdsF
WlK1dK2S0fqPcxlfkdWLO4+4sTHHMHVru7lTfWdk3s2koisnoioz2ugK/mSNPT0dAad45SJIV8fW
TACYAOphGV8U3Bzw7olOfZUfeSmdNjPXyV7IQMw0+uFjb7v/CXD0g0HXEtCWAbZOHHuLyfi3vgkO
zXdf8t/qtaVn/0LLUF6AKxCmRzW8E5f/DWLUiucbWFj7GRC42bCz1XxSuMlaU1ByHnAsSBQXN2Y3
eCyzAZRd+ezatsIxgy3W6LleK6LSL7QB39PK0Jy6JS9iFrCnDJRY29QBAqKF+ASXhqAbAKPgj9AB
KUqcr1/ueq0Xqeeq+K5g8T5EH06NN5q/hzZE0DN8LyCHYzelb4KZfqMQbJVQdlkh1eIoFWhMkAYi
NVWzKSu7aX+FgV2RYjnpSiZd+o8+ncGR0zIYh6gjFC4NwCPs5kF1p2iz/eOtUBmUy0m9FYCJd/58
Qn/Jz+rTephgXB2zNXGhkxoHhw3KJAaYMIBp2O8IGrkmxqv02VuhHdGvn7xQTJu6O6eG1U8bIiDC
Uk16ddnVcCEbxm40pKu/shtAxHjheeZlCU9+f86hL0rV58J7FH1/txogIrIMmDuzOwF33u0OOnSD
hsMKu1nGwjtQkaS/2sLOVHfUhu5VOUpVMQbE4jEVTggb2HnqmvjaRXhAIqkxCKf2K5VajFC/+r2M
GsXSPfBazO5afASb6iwtKXsuzPKvDPQntYhbuLfPKu5t9p1GzZjLNkpP0fLs+/GTNeUtFv+v5xmj
icphCJSM4ve1v8XmO8Yj/8jO6kUsz0/bXvwdr49ryJ4redLyAWYvCaoI+T1AohpEKLtgyfHG7PQk
F5HK35ntEFMAQ1AsoUs5dhXvT8+/uJLPFCI3hK6lb5j1PzcpbCEiIbOvuVSsKVg9lUDlmXlG7lkk
Rzu3GH/8JXAnEv3OsjbJmzCoIqVTwNGuPDb9mUyl9qJyEGBQKl3KF81gBqxaWnn86ZQiFUSYPlE5
Vtvpwon1KP3LGJRtv/xfzJJeWnZEFRz3p+Gn4r7t2S40jjNAB900wT/PWMTuMr4iWjTj5uTE+ObD
aHrnQe6tjdRBqLwxkoobyaXOITYKysvC8dvaGaFBph2Muvv9P/9a/Up20M2WKnlhzpCG+j+AaE4O
URPri0EfKlrkxmzzCtVkMh87bre7BPI4WMmb/+ztmpRPJTEtN/llDBiT3TpeUBG/UKjPRML+gbtU
3++n26nEn5A3j+jQk++9VBkLCSzpZa9py9Pl572Z+0bVwa6IAXHU0iyxaAjqZLYTqHgSEv8FG16q
aB/oM0vceqZIC2ZxHgyW5Sd75MGheidXFQlnvXtRoLAlgruq9LPSALLJPm/ooc0ojfyv9uN3n6zO
SBqnI6ZUI6+dbYu2bDNQD5HFOdW9apXTkJa2zfMtp3DD/0v01bypfyqsYHQY4K9tZlybPY8o6ur/
JEeFEY7oSAGHM9d8TdB3idIhuKeNq53tCmmQbUv/DYb5NmMhvQPEbwtPZDmSR4MOBxdVuAP2kzcu
D19IKwu7BBuMPA4Gp2KoWOYHHrW05PdYozlDxRinvCM94Uz5G92E5f1ClBt2lTbex4AFffCs5Gvk
JU7nXm5eWbgAykrup+35WXnpwgM8iPYl5+eS5ZRyfJSj5vLuUKUvrndfR29AQRsFOK3x1hhfhxXt
25t0H/HSrfgsEFNkEicKgh6cTpxQczOvP10Zubk7SBxi93KX2vfh4tS4iPNqWmXkgbMP6gtAPe9N
+R7r3KUAori76Eie+JwicQJ52abwkpZVNyDWET+DsV3hEdSgOpfp3j9MYm+koEZ5CbF5NKvhu/fD
nmAXRWTR5QnV9bOEvwTxR7q3XioxkJXhpR8fL+R4Uk8YVWuTJYo7qU1dTB3Dmx0GZVjw8FvsaVCR
mcNfeDu1RK9eMNOlRHoDXchif38zNJF2vhJXiI0HoUChqTPClZ7dJVzP0GvNUpSuI0NZoMYrjHnB
jD9qC6z2lKX9nlfx55VeTCRabhni39X67XKNchFDaVzeaAtGY7USPpzDPaYU0ZNMXjmsWnnkLTp7
mtu/cWlGTn2wcRlXItSuLLEgIepolpzSxyBaf4L+maAky3rlN2Abe6r3cKaT+fFL71yjBWm3oM1E
7UQk7NeWjoqeuvutkepozyrKspYVfBbvJoksbFznzXqmgOHksf8spC00/tjuDCGDkxddkgPeCb6M
7UPNi8d4c97+Oy14kQ+HMGUue1hDQil3sstUBhtMDHkq9QTlRX7AOvpRV9GPKgWo6o8jiW03a9P/
jGxgiO8W3qja5jzv2xfd+fecSwu5P9eJGdVGZAn1VlucSz7u4KyMpYWH8dcHUymvHr/yR0fVmAdI
Xq7R+VHeQV9N0TprKZO997unguOk5hs5gtT+F1unq2DK5Y13RSNdxyW8Ij4u9PgGuy/8qF8EU0b+
5/EiWvRI8Dp8oG86rrVrWovzakY7SfKW3LKvdGjn4pgiYacsJq86tpgY53unYXAm3SFzPTtoXAwT
I8fZsT1Ps1gO1WL3xUsCsPBRVa8C6bBGmQgcFYFNtuyleDI+1FASIxZytxX+5XPdSun1ZpLhXKxP
wMocxB2xCRF/pn/xQm/NE6xqkhdKJUcGQ6VzSV04fYQK3/vH48wfeysc4T+SVQD4PPKfDUkEasiA
OiJXpmhQjV42LHc15LnV4aitkn4HmD4fD+EqHlE/H6uB3hmutuD63jBByusMUqk2uQDXCm7n7EQS
48VFykbVyED+3YpYNbEvE5docV97HgsjLrHYcanwQt2lgfBPpv7ludkIcRL71MrTJPGq/gQAIp+9
88eGuJPn4wTisudGWXqEJ10A1/XUbFp36x8CdFxHdXhKeYnLlv0qKwUm9d5VrjV2fpEZDV320SZO
ICciiDzI/6SN4zk/HLivJwnOLxbkRwgAuNZ0OCrMLnf7ArSqHgMWle4osLdarsWkrtnvWvt/4Ald
QjV+tyemX9gqb/OeQ0rUBDhK/b6gjbukFqnokM2yUDF67Own4260g4vCN13OZIdEu5c6fcAaVNmk
iomWnryYfFJhd6XMLtM1Q6difKVn0ZmxCCnBM/tKkEFPaITylypxbqqO6/bukeNjQwGWWoF+YeEm
hBwHlQHJxE6ciLxl8YDmWzZOVgBhVj5nFmdddsf0X4oMIy6h2QStdYMj6jWUlfwIrYLXKbOp0bA7
WMjCWyJotim7A7wwoFMRDvYVG5jFh2y5gz6+liu9chiCKuv3biA4sOQ9e9NBS1My9BxV7EU6cUeH
wRT4I2mNK7LKtsMBgofVWPk2ygsuCiKZ1rCY0w/cqH37hp4MOGx2tGSDB/leltjHmVdHAzYkxYxL
VvEBkinXUdgcYMdDOop7QepuqZtJd6+l+fQaihXkRKa7PY3jwY5AoxYlYY4Dj1lw2KZmwQ2rYhQ7
IkPlMP9Hl349pR8BjyFjT/YJkYiVi+wUzOK2bmIfrsrM+Klv+Z9GJcOe4fgCxQrd1CA6gJym1H9p
o0gxyMV1Cyp8IXUjPGEKknszt5Z1duP0zlQ6dYiGfzuyZWu2+Ko6YO0gD1cSE6AXX16mFCFBdBHJ
Raxgewnk9yzIzoyL2m24ih9wC4S0A6ES6zwQWJVpQY6EcxmZpLnHKIgSHPg+8E4oIwy04NbbIEdW
0EU+1Qi8E6aaB7luSbY9fyUnghDF9Nd0cyd/fcI41+r+JXz6i36afMiL5G/ortUZovYmtzG0TAn6
Coa5qvqJpeqClBpRkTHOi4g1scpSTEUrhGHT8Ct3X11B5i2Au1B0JATt471wAgzD+oX+pt2jMZFq
sKe4KsrJNZf4TB+zKM5/Rzdt73tl8432anxLp+14pabsCBp/MvJ+HvIdUKZ94UCV3YCMHUh+lkvB
WvECKfYGFj4O05zOS3xSg4lBJZAS4cEWCJEEEvQ9oxOeBvL2ZLlyVj64lsgZws3f1N7xsixFcC5v
QFGRxQnK1xKrU5en4u1K4likYDWCJtCMCsB5IujTK9aZPKNlf7E7hEKJ9mApnef+32JjNQ1WL08T
3AW6DasOo/Ln3opw5ylgymW7ObFi9JAuEr7m/lzwGfFi2yAUfUYze/hz2PqdYYkaxZ+YjyRiFFNi
+0E/CWHLMYw3DyIKfC6Sbtge+4scK/8S7hJj79fniF8gXCtjdLYnyEKK4fEMaDh7i1yNjsjCWYJ4
APKjC27a3xtxY5fU/oe2BDa1XZ7uoRcyJiR3AqcO4La1maZ8Y9zODDti90/kWAKg/iYuUu5JapWd
rxlU4IDnzJaEN/Ep4uImRkay+nqZd9Mywrkd4YdvhDm4MQsh2Df1s930Ed1N0ARXvaI+dyifArh6
X4RXGLR39BSd0+hxXOlBW3WWfAw9AnVH98PKjYue2dpalh/v/VDFX1PwUOeG1koxZiXgwqA853Qt
eD76gDRcA3NgDMkS4wCBkC8RenrOtKK7Uil+6wndHQO5TZ28jODg/ihzp5DZczVRFr5ss8k00Cp/
XbBxlYK5tkg7iSxCcguqWjGIh6yLv+8O6keE+SQoxxwf73EIPin/lcQ5VN0pYKd3ngpXPBsF8Rxe
WC4kz3RN8RK19qGHMu8NKRZP2QadnFBGcAS3LW/1Pkz2710u0QwPXbJb2CL+VrCZ1fyK9XA5kevo
Yq+JEMmgy8daL38BzOJsNlKNTbqjBY/lqyjmohYTjGhAj+Yfwe/QQ0xS3q42LOP8mTovDqO0YxDx
qYSsBWAHsn+Zj9soW5K/UCl3axa0SaJgK+LfPX8Ssx4xODJpYro/pTZuBZuqzMHkibigC+NrRhdO
0yJYSVHPAqnStRRejZ6vg0lROVnght+8pmTg8C+3/jUzJ8KxCw08NS82enDWzUUeRHcbYhsV76Vq
tMX5sKI5U0cpprHuJU8sS2vjCySBAfonIAI6XkBzV4f/FjyhVNghJfnjiZxHkQmlqbRlpERulC4s
wLppqhu1i0LEihE53Iv+6Fk6HPuGeaIwi6C/LopgG9l6hNheFeO8xu7kfs7hTidb2h2HqGjxjlBl
wH0XQF130ZvBjjHd6JDFkMGkChwx032kkS5FT9tc4BWLhLZiSYcKqg7B7u4O5P0zsDdjimLy+5jC
IaWW35pHwMz5q9VK+B42SwSZDcVcOMQ1mGXnc52+gOrtJLWCLIzW/suzFbAUTH9WmzP7E+EbVmzb
eTWVNwe67XPN/f0JxUwTENkkTFne4YC0ozHiwb4hfTsIxNyZkOzFejAPiNrgoE4WhRrPpakKvF8j
Lj7ub+FLUVUARXirICAFC+jrk6ChSzZJqCtjlzB1S3fx/0UjIwqbhWDu0eO79N5TUBJlZD/LEHyL
c6jErrD+JhTjpKAm6Xc3q2aFqSJWNObS+gcy7+zY8biIOMhMD5wu20ku13K7orkDA993y08XJoRx
cKeCJZB0s2sb4IqEo/BDcSoyRedcVUe9Az/4UA0sUv8hgIXkkkecgvOWfiBVj4UZ+hhtGlC0CfP/
klnnbw+5evM2+PfzkTqDYIixC5NSqUxlrkmmVf7z7qqLqQvHOWj1nuTRu0hjALHHqPAJtXgiWEZY
RRTUvmtVbY+NEVFWfGyirj0K3d2ooZlepjZaxPwwDJrqCGPRyldeUg6Kr/MKrSHUzu3stPb47sb5
SFV9E4dnR4UpwjF+di4FhX/YBSRCpSkmglluH/lJvRpVOKWQ4lR55XzznHuZTGC/WBeF96P4J5va
CYowkGdqx+sl7Q2LfUoDiOH2qOS+eCNcGdbe50XqUxImukRGT3H6vpgz+tOs/TfX7B5K3bLiz/KH
YPRM2J4RX5wsSd8/ZDmzxQ2y6KXxHLvxmKX4Ab7aMT7U7VafzvMoJgN4Ty+hETwxBSHKzvJg0NIS
YfnkR/Gop4Wr8mweZ44waLlk9rh6Su4kKIEk9r8UUCKFFSKEMEkDLtQAbe32j6vS8dLWDB7j0+TE
GXzB/oXloEXgXnR6zzB4MZzfz+Jgq2gSyjHjY7ZXrA/oSRGlcJBebL7Q+kJ27cD/FvTg8wRD7VyO
IevrQL7L7frEUAuWGxs8cuPkY66FxnIlPW2CheWBgWX3OFAYNFBTdHjVNHn9yc7RAW2Dt0dW8nqQ
0Yra0uk/TiFiSki+iAiYZoVUdzBA79mtDRXIP82E+dCRevdVff1EVk8MMUBapMKOXzPWYOfpEC60
/NP6ZvI9/NLqnPez3QCj/3GNy9T1qhJlSSr7i0EREGSEDxkDkVVac7Z6Xenjs4/NRNMEdRsyqjwj
fQV2GIOZk8lSkLOE7y0L1mNJtEfo1PH0RNWWvudeVuXcxBSADhqdVSnC0+ywhLjrJ968TOXKQfBn
3SM668Fthlb/RWkVSmOrz5r4UpNSknlctXaxw5gb+D6+ftGZbIVarHDd6iC6bGdTTVqUoSfvl6e+
4sLofDXS8SFi484RpsT7WjMsSXMcWW/pYINTEKyQlPbfchZSmT/ijwkkT16ypaF3FGdvJY9Q/h4V
OPTy9c2c3fR/P5MFYkNHRKJNrnuT3eAJ57d/PErODSGDjO83S9Xv9wFTONI5OEGxRyf3Dgd8nqss
lIVoPU08F9ZEaBRkvqVWNj1VHhGEGMS+Kruaz/94j+G0aEDkpmoiwk3cQQV9MCbjQQCjtRi6eERV
Bo0tFEc54mO3Z4RbO/pxiGFRyg/m5uxwWExzbfe5+dvVqoh/22x8anbFNUJU3s7BKMUgII1gam1X
E8TOsPOI9Y4bf1qk7hKgVXb/VsqVSxJbbDy2g9qvNwmGc6i7T5e7a7F1snVencmciLrVyKoH+wly
2Mwjnaq9h67XVkaIjIoRv5Qswx8R0VsUD7RMO4SwfzPO6z7JG1GGTQxD9wxGqDs3mOmWqaacPwwB
10x9z5ZRatSvy4nRABLiI/X9JV0wvp/r+9Bu2ZesfOyK1e6/VGmq+tzmmIk2XYhIRNu3otsMwvsq
nBM9hVhpuptiKBBeXOtM8dsyULTcui4br0HXzwjRfWE+KHeJgew1KP51WjkGg3cWT13b8fNKKH5c
F6LlXKdsuj90sS6RHj3rwpZnLoH97ruyhJzwxKC7zSSmtyKH8o6Sp3G2qSZYddi5GOyDitWZfW1O
dmCx8U7Qowvj4aLKhquz4SMb5J63mfMqVaOzQslrWyRu/wfdv/Zqg5p5FGfRdABa0SDpSAWL/8Yx
JuKoePOEr8eTeQA0ZzxQPWRxRBs5QA7FFJpBcy+ss79BN10rxy5uVKK8YqsMLn9MnmvN4smf7+rX
wVNyR+oYTo8wpBI0rzq5GQYLB48ew/0f7yzrwfpkQsAR0i+RAPU4BhqDHup4yZ/AyHhUASVEkBxk
HW4DaWjU/MhT5YyKIUD7ROJTXHvlv6r5exhZyGgzNaf8FRBwdle3wRMe68YBXVZmjHTvIBAXY1Do
AQ1VjenvepUVuB2UZ1NXmjDRE6KdvQuOLe5wy4FhhAIh5iq6y+7WCNBto2PlkA7kZrKrpL8CFUxz
NVDBCNcjvyqfnrr18pc3Fmxhqo9jSR1VrVXR8Qm23DoO9pFyvowEXrkXFjrfOQ5CXFEAFgGfgp/f
212Oy8wMqxfzgDAUx+H+XXw/vWXOBtz1Uc2VdkvLnFV/xNTCL/W7AK6wKKnvZAyDThinBD1mUyEk
QwlOSi5daEeRt/swqAt81zSa0gEproGMneVNjDn+Q0IrsWQB0DdqX3GIBfr89pF5tzQYeic3fpwJ
62/g+OdIpyQNK2Gtowli9rwTk3z3yofUUcBzIMctVclGlRn5pAaQUfie1zmClnUnUV6aDUQK/uld
afmZzybXKqJayM/yLgnbkBI/d1yNcKBKAqBVdU3UU3sUxkdH85eNk/XU+x+J8WdCIENV0t/Lm5bK
RjykcLN1w+lKWCoZsHZvB4zwR1keskqYMBt/eyVHzhxPSdsytPbcYrZPtpgsG2PzMXjpEmRbH+fV
HUQzVe62RD7eOK4R+rRVO/yznlLYWlAykNe0UI/tC/ffyH+bGWW/8tuER0YqqJO96Za8BXyAdPIX
lwRukwF+6YDJFirgpxH7qHnimxBz8uA9+bK/abPG9j4CQtltfErcE5gIQuUoCm4+tvJtaxW47Z8t
1WwHhzgtfkbZInUieyIpJMWpT4Z7Qk5wKK6kjWaNwnfGNMuVGES3CZJev0Ltd6+OR8wxPheCO9Yt
MxF8gY1bsvdur+rkmCqikxnFKOLvrAYlrIx+usCZXKiVuofSEBgMykEh6jQA6fUL6ibMxVNNlnCE
9Fs/qnMUhM27/Dh+pIs1KEyCEcUY+IYJpesqNIs2mQTo2m/r+Qh23nwo5EsrNZiZ9552o4/ttwUW
prrgiMMgJEisfGTYPx2sZJ/BGD4KguGJSVr60TxwhFmAJyVWXAjMRNkCmdeoyqH7M/gi+bKqBGJZ
6+ME1VZ2VoZ4XqE0zjprca97Ki/tdMTG3M2odT05LQJAJ6hCLF8lqq5n3urh0MlkLKFb3Lc+7wrn
weve/CaBJPqVDZgQhHrzBTlUceJSHlsTMfG/4LF0EFJUgKvnZnh2cn2Bly2tJ0RPRvwj4pqsylja
iTu9lPLFs+67l2Ufwd0CyvwyOGz8oCYVOJgao3waKgcnKpMrQcrFBCDnTIRXKBIynoh6lKboL/jE
tHQ+gBmJk+SQJsNggHtnQ12n/MVUx+a3dwYXnXh4M6fh0OLmb/RbK5elE0PEYNC21MGrvpRtv6u1
paj2G/drSYWbdohF2KwiRLOJYejvHKiiAjjL4Zr0IYBFBKtki+9Q8NoMVxHW4vty6uF5adx4HnNO
imPGp7bIdRie1ieu97nWKVOjf7MRNqX3fJrFkrhe9pbIje78Ydt+4oraJikb7xcohn49/x+ecjSr
+gonxUw2OS/TpTPOMjfdobCgcYVutilnFxzpsctT2HutYVPOOlLYkinvc8+Mxlyn69auSXbJfN7y
aDRVIfSw/pI4OKRWsW7ISSsce5tZ1LXfI8F0xKdCUgzGXAMvRRPoq9sSTCwHBcu0stLHenSQ5M6R
2/bOUMdG+PSekLOqxkdRrh+DareqcYIxMTb+Nd+IygZnNmCZiM6xlGF0dZvJtFbc61XrY2WxzCzG
OjnNNqqdubaji0M4NB13Egy12s4bm2DiDR5SiF5+xYLVhmfPxnSmxUgRaE0tJDYB8eh1UyD5zOjD
G+9bK3bjNBE1m+svbA3pIXUW6OmbJM4oJVT6p0MJqetB1xJ30FGSzJ88eFIvmcsBFfCwcJm3cJRz
/Kbq+ddb5uE+8/vpLkqBU4l/LQ3bXzlHX5qv7n0xbA7Ao7ZomJdXyy7s7yzS+lrxoFU6VV+QFWkG
/UxcwSW5ceK8fYvEuLdQxKJSKhmyBsrLPQlM73gMdQwure5zh9IhKGcuMjttmp3FAbW90AYXRldn
HiFW4XTf2bJwshwRB2+G4Go3blaKmuyR3KIYO5Zw1hvOUR5/UfSn00hs0IEaLj4U9t35Ogg//set
UEeHWm9l+JBKN6Vwr896eGv11CKJXIfHKL3Wwv4Yial9tWepS26P9b0SafQxfJ+p84yeb5buQyX+
A+ZYLwnSo2pNlkkwWihb++4iiFRs0IvQs0g1yzy8HmdVRpFy4VsGjN5UJl4jJFdv6E0jr8rwc09J
GkQNgGTsliUjyuJfvW1lhxRBr5P+7PMuGqNG6ivNwAZoSXOqohAb8xoavwUgpWUqsFzMZctUHcQS
D4cT/6WzRcbtrFc9Ha6HkuwqvVGTrzqToN+uRCQQxzlOuqq+rnTMvMFCuDQnIYaWaFhlaiv9f6rU
fW4zP3ZES/Eu4T/pxQmVoiVq1KZriYbm0ZXPwoAQU1eDNkZj4AeKnwodijGnp7XIqyf2EOH4tChA
lIP0HFnVphIBfWKSRAvGx7o2Cn8ysZtmM2Z4M9TL9A4VYg5kbNta2kwhDT2xMuyI+FT3mDuZHLi7
e3WoZSf1ebxNPAuCyByGr/VHJqOIcNAejrUrMYkdXnG5dPY4NyS4XujMLLtSzWvz2KTgMcxr0lRR
odh0pyCVbNr7OXqvkTV5i5FgBa+QOPtYu6OwrrWUD8q8SfUc83JFGU/F5oeOJ1hn3nFf93BMlCgK
5V8EV62rkDVaxOIG/XID1p2N+7daqig/jSC8SJDVKNic1UaK1TGSS4LM8RzHWTjl+B4c17y3gxnE
MEeEMoA//ix9OecWOty52e5EjUItrfNXWqwe3E2Dn4bMLlOIk4JkYdNMG6dpGrV0pPG4gmCDbdfS
yyHS/fqZGDCTVIo5Rc6acr/vWWguL64JVbOVBUKeIQgqHkszCmHlo+Uujuy7adHXkFR1Ej482TpL
mkMGGk7wTrcKBUeYcJNT4kpZ7NPAprUonMRmR2XpzL9vIod06TQZsoWKYQadFIs0S3wYw3NKGglz
HuRz26v46xIU5Yqj/1+aArJySAhobcmFhKyXJmt/4LEBRlkN5/gH5lv11qVDbds4W8lcECMg/uWT
FcIPGPHrrfcgUnsJqw+ZuM+/OrSCLvYeOH7P7+xD8Acqwh2SzO6hwJ6SPEeJ9blyawKnl/t/giLQ
/IAah2Fuw6bJbcEGaQuNNAmr9De5AQORbDuY/i0nYENbFTjVD+MWIL0WQ/QQ9bWjtnjWDSxtwtDm
Vciz66R9ZNWLL9JGus1r90d1EOJNrnfbMTq8xiGKnF6OtZ53+G6Wre+DZ/5qwm3rklA19cnMx0cM
meY57VJgWki4ET9DaAGm0ulHs7sDwi0SsMCrSBmG/STAB4NFBSKqPcLA2MOA9lXS7zebxbFUU72j
X88KgWmDoairQ7CnPGV7qIc5V1gvL22t1v9XpNP21keoLn7oxSpD6y8uZV/DrSvgr/LMsC7+Nqet
/bEAx1ORUs+oVM7xwpS7uhnXHZpJhqNm5TnYgMi1W3TeKhgbBJJLiLVh5j6bhuz2WI1H39VBibTw
Y3Yz7FKsXuJrUPwPhjvWO7ZcPEwKT+F7pbGnLtaOdol8zsMkL0xplwpLz7HUuCgape1WoyMu3s3f
2pbGNG/PiuMhp/gqiA0P3TUkIUX1xmjiaqUEn9oDA7lQgNhd/hmzoyicjtq+JwL9JwqY6tT+JmfG
eJ6OhIfIKUxk1QydHP3/tmKKdO3jHjucC8oEtB2eR9+ZDemWK0EEk/i21htS5HR31QiGuYtfEIfA
NhPAU2r9zR0+tFyhWZ5aQphx7WnUVjLS0ncrhtgqSYzUIGzsLH6j/tL+E8kno2lr5ukyT7nUiSX3
wXkcznccvGP3nOkx5JbjFvfYXmS9tvg82eVSsw62/C9QBPXb3AYaeqE+1Dmq/GHTTNrKImjZhGTA
nOJEL1EjgFWShGEjCr5zqnAk4H1VyqxLhX71r3fnEngrM5CWGswjvGDWo3dOsqaAXbiy6q1HPdt6
URZudmdZTnLaZSOAtvxMuJIruL9Y2UYF3ePvDMDJwVJ118tF+yhXZie9n75cODgI+y1IfsFaOL7R
/E0bS4N8E4FpElugz9Om68Psc6ySTiO+rN6SR66a71nCWKN021LZgN7L/e4BlB1UjmShbzZnFaNC
N53FxQjeOuJQOP60zi2WkNmbVVSZdW8tCoInhx2eG1+TkI+IHWK3bV9dx8MROGVDRcQtVoU9xtQR
hOSzuwYPwNK7uExGaRoqGxl9mjrX/MF0TmaAqgoCpyq1wvM8o/79IM9MojoTTZVmUU+kLseiZBib
8Q5uD1QAGQtLq89kK8sy3lVGlXGj9kI3hj0ECEkSqeZM/R/BbxQ58WmF+mPeNthlohfvJrMJ9MC5
oUhGQIhZjmd3aWBZNip3RZDyB8PAmBMYRi1C0ME+dkxZVqn58J7dDXM3553aw6TDrtGmBXSV1C+R
ocjeg2YKiP3dwoTUKoiThLMWV2NgdeiVZ5Zyjxy5QrwnxQzXKLmOUx2gms9FYcdr/rWR5tvjNrW8
AAgOgC4CJ+Ei3Vt1bjY94J8HX58jHRU0cXnoz9nAga8xW0VC/Onu2+ftqSWCIjPzyuMRZG2fl3nn
9v1c498xXhcZ1qK1b1vF/rV96P+bTw943hXYR29OTJlx1iezKonnrw9qdM+XutX93YEi6zhkuDal
NMfK6xznEFsYP3bNcAMzN6dB/M5MkqKpOuxyb+ZAq/j3tWrkrbDVzTj6+GcWIVFc3QfeoL7K19dN
w836dGFj2rY5yUcnFxA8dyqGHMNiIOPrGExdjmy1yXAbeQcdiLx5RIvKr8d+VbQJamzvMuFsu71k
g8aLSqO+F7w6gDbjbU5jqgTCvJl4zNQZT6k+EgfVA+nlcahlPpVtIPSDIn0fEGws1yubRdgkgwLe
40W5FXedGgk2d6YCYk37yFAhNo8h76GNYg/oRrTmmztNyn0N7GQSIA13pxwcdKVj8OfGJnp4hLat
vMrRSWzMyM4e+KAVOj8PP3bHgu1zZp0bAJcK9fsHTuHuUpasMZ8b559VBjHFr4wg0v7IFXWHcyLU
s92isClNZNhBX4QREm9a15X7Ceb3n+r/JEvmBJsHBPvhiwt3kytVDv+q130YoZrvt2U/daRZj3tK
a2hAryJnIMh5fRmsq0+wHtT3JARkcG61xOLt+G2r4KppPo0W9jxH/iP/lz1OjVI4iJ0PX2T2rARQ
b2R8Zm3OjOGOAo/UZLVYI/mlWMiKyx7C0OA4REH9hn52Kv3k0ldxf5kkNb7WUdHlql7v7irbaJC5
3lmaqyadb7CtIjj1OHHhYda2wrFef/r7HX18iix5Erx+BPKb4PeGl1n0uwFxx62Hr+91BFNwIb4H
IUUBLI8HTkVg2+oItgulizZ4mvC9cccAFJTPs9dpEK4xpOojnfgzwtH6ZkyXwye3JM0wYE/ahg19
CPPLkJBmPDEZeCPivsbgl3pjskF62PlmxgggA84ZlMtXZoS8sIH4zDprdghfQ2wEgtjMJcnyQOrf
9vs2vD4zIUt1itjuysDxs0PzkHsRjPT/l+jJe7Z5ShbQJct8mWA0+OqQqFjdQ7Ilb74b1Ub5ARMr
ciHEuaoHwsiqcQ0612Q2/NesprBE/qKCqiL+vPLacXU4UsOs2B7Y54EVCE6wsGUH8c2xIZHXSFh9
ERRZoWdCPT7l3wxnd7urNqABjFYmnmIth7wabQPC3eTm672o4zP5p5hQ/6JbARBqieRt8o7BTgSX
gCv6YIIvpAnU+1foT3Uy+vZnVQCdwbC3CFNftS9x9806EeM/ZdvoQgYJrrjyGrOgaNbtYtjys/5M
4E68NQjjkWCVnjOAnZym4ro0cNJLJKWe7rJWlIKGhpn0y405pb2V/gVDVQ+TyVOFoN4QEB56/mdh
gm4VvjeLfItuVw+ET6w+ra8TzWtIWfvY+DHZINR/RDTGm/KnV3YPIazPtpDjdmQ5MbdLnmg8iYv2
TtIsv4DqouZK1ksNjFgB/+6Z4VweS1Y0JwBjbXuPy2xci1GE/M2E1KteZgKORl2PcmUNpgINTpP7
DG97muXBpa69VFfCfnT+7TnNG205mgFT7okeOnpSPiU5msNyNsOlM/7Yi/OLQLeoE1lg1QARohdV
j2k8IHt/EtktiUtkZq4otw+scfGgPczNWZRlr/M9hSy207utlUM+Hh3w1WnfW5Hm+QnfNrLjTkrd
nS4uZLh3GX8wMGQ5K1wiChmZRxkCamF4ejgFGqb/NqJNAV5fpRHU9TDa/woBCMv7/4dlUA8ihEeF
OJTacZrd7D/q+XFio3qD0j9FlkV5T8rP7PaIvwfzdqO4MRWLdP606JLIXU9yk+zJJ3VWrN/Dty3e
XpILn933+Y6y/njGJv9sDD+uxsl/bFNh/3tWHB8ddDacYgduyKi0U37Rb6AjcLW3K9+kmES5gYHD
khwvzDWxdHtvG7IncRVAD5la6WbmJ2FSGAxJ359GCGjVxpTOuOXS2trva2hZ3cIzPTxutEhXgixm
OAtvcqRj4dkZky2tMX70DfPk9fbkhOULndb6zoBA9IZYsMdQfXZsnMrWDkvPUwHC7uizRbGdhCc0
3FUOXg4EsFoCFen3dMaG5ziE+iLN86KJpdeJ6TFovbid1HM9C2tdsnRT1BurjQ//ibuHTuIT2i5e
HEXanK5Ab4VX4VRgRT1s4RzXeD1QPlobUFtfHSYKMPeAZaA83h6OBkdgnUQ+28L+9hb65+2duhP9
RWYPJ22uacPG93CkiDa8/96M5JaV4gcMNbaXqE+7ZGpt6LPFOx1CP90f0J9RAa2qW6ZZkKOdhsMl
+eSC4weaiOF1o60sEj+EbyH9c+7Tg7agtNAGSLO1ck8FOnAiTZKOU9/LRhXJjD7FL3K5csSFbe2v
tF/aT146JS1gDJUJTpdywMarhYiFtavJm4TH6ngvNYxFmSp6yuMSGAwoByydC9T5yNgrkUEAaMU9
oowdUrucDfAZjeZ0XRg3m+TBygGAs/OJ008pWZTF1tmt9CQI453zaK+qE7DfX2TiOO6CY6LXdHkJ
/L3OSFHf4rKEUFGt08TbiG6sXal3y84LeuaRrSri36taPJGjzXUlfdLzoroyG/LWQhN4RzHjmsi9
SvkJ583PfbJnz7/x2k+7AZh5aEHxQ4lJnOQbGqpksVsxlXa1p8233vspcNywdDlSycWt4RiLiLsp
B1ZffbnRrm7EehTLd7e1NrpAmc9sIRjVlSOpAeAxNPIGqUePfuszE80I+HW6MH/q6GH9VGYkc1uO
UFGqw1ds2CxmQDYmCNwXC4gchSTpi8UNg33wFuwmWrmN5QYLsEwjjzw/XJLq8lfzIniCAAOUwwg1
qMb1QyJQTnmLfBFJts0uAf3x3RU9qgKSAVJ1XlHPoMLFrYVKX0PzN9xy/EDgzUiAinjfTZ1ZAj9I
Zt0aH8gaQLPGsdXsiYQUuHNG4lGsU9C2lDWd66u64k0Pbk7QiM4t5HdEuX9Q/5ZezCfsqa9u/PUQ
X9927gphsvxvOUfOcW9OJ9XhfMZuUpbuNXGER82gEH7PqRlOmn3lWCXj4jLI6NHL/FOaiaixdRB8
GZoK+p69svaHLCJhvv/raGt1kAj7rXROP7VFXYiSdN2+LHu2Heu0UuJUVAvmaKRqi7voCydGx5jd
9JhEuZv/1fbSj5soZKNUpslczORVdx8PfUSqbnO6Idie2KSxXzKAraqi071x9R/PcYF8lb47FGqR
y9JV/kG6MbrFb5r7+d+EccLClKNvfwm15LY70qqxDy70ArNEZGP88odYRjutqDe/GPomsKjfAd73
b5KATclNKuyJhPLIwD30z0aBHGSecKrL/Y7I1aWfkeYlYjgeUkDc9Nozjd6aEkv6l2+58elPpnxM
0CFCul80q5q4KvyTJnT+P2oBmen7GzbQm4BWp51ngpXMVpF04IkU0chnmGszT6YGxy+wXDFJecqh
XWs3Zeh759hh+byDb+vHbugFYrT+IIfTEiGlo14X85hlZ6NJdsK2N8Txlo+eENLZLXW09J1quEFc
JVqzkQd7F2D3j/a7tMuPh1bkga/gKrnTIDDX4CZD48tONXzyTXMP1ge7qQdrcopp00/jwfmj58e0
b3wYPT4rOtc9ioChhV7PzzXtuSWrcRbMv/5duEsg+ZiXpP/TmGur+ZNoNY/B4/4y3m/+NnhD5+9p
NdAhbJ9ROqpdy1tHUxE8rfJa2ABp8Fa93KznfJLddcepX1IErtMm2f2SjYJ98KHYh2NIyK5hyQwT
RAonSpWGIFmj3d83Q5PbYWvP26xLJ4Uytvc7+qku81G8MxtFl0EBcrIpg4HTj/H67TcvPq4UZ3of
Z1taAPLVAqyZt50EGpPd9VwAkhlfYISQomF8pIJPwIU3lT6E/aE0bvbLsf3RfrHTkmnGnQWjFN9k
PYwUi2wUmzqHucwPNX5hvcWSws3N2KnFdPFWhm985v1OYwHQ9fhW1hR8wjnFixYRDiW47uRpR/yS
Ix8yMnzgj6DrQGNaPq32/UM3XpUFQjW+hZK8App7Rydk70qW3MHh6VGl2VD/7ojL3resAJn0Khmc
76FLtv9q4TsBwR+/gGqLscWiGX2/JMtvbFI0jMSoisC0yyTwMQb2sElO8V2/kA98RD0LfGHqlMpu
RIn0l6SlLD5ePn6aMTDGwO3j0ib25jI5yvX6p2FflyfGBRBxsCVMxxzWSW/gOXrtF2FFKeFnAkJD
No1PzIOF7h0PQ1+NGujNOI21UqBytdv/Q80Bv7Rr6QUi0skLzFlc9jt3X51l4Hz6JoHkhp4cdO3O
5ecrK8xm015Iwic4s1b+AhdSDYt8V8XxuqEc58QLjN0WprEw57ALwJaMKKpHfpUER7EmUrfjM9hz
2J5DOhFI8RyVWtgX+02ji1XTR4YWBFLT86/wa5KjPPvzuqTnpaEI1TKvJgbpzBl/EKd3aGkkqSLg
P5H7mTFDMQ1/LQg067ZjaGacnrz4h54doq2TEWzN4NRz9OK7/4uzdd8yQrJ2prZuYsotet4Urw4u
/dxq8VDftcjifaJQDe8WyuqX6/3Ub9lv5ew5ITTAaV5jrkvugIiZmSqYV5BLY6vUW6vpKZY6XHob
W9SHrly7PLniWXFy2GDz14qJu8Qi0FvAkWA0/SLgVOzlM19/YdRsGmEFv7uioZCVIGXiBQM6d9q4
FswxTp4kSjTogiBh00pSf+kWjm9jOErGuelGwaZjQ2xklbq7UAL25Ls7p/Iyq/PJn0u12NCmmVrE
anebmZ9MWS16DnUqkB1OW3i79TtDC3HO4eaHGQUiOnIzdYwWf6T3JJWG/xboNTS8e1ygfNGw5eel
VLk/75iLjbZGSAMZ59WNJGkDRsuDf1xcbA5q+797XzXgKbHNqLP6qtEmuELyQTolKirUPdbUo7tM
bCVbMc9zF7GroNKQWLEMkQL4OSfeD4VzY75/PnTfMMbrbtoVBNCrS2NyCDPFM6RL/LaxMt3xyj02
+Nz5kqikZi69tuzw/3Py5uIIA/I2Jr+bdmw66ndqPFaVtP9trPQK7FZarYUX6b9u8+TDdb3j8GgQ
bje7I5Ws4Du9zHyUN1m+Imf8gMyudOm6J2wjnUWl6ZGjXSRYO4GDIIiUz2A+g5rvFeahH55ftt91
URp3xkX/69WvIVcNEIiEvwbLPz4M+P57aSVWa/lz3oSQB/o1sEvE6I2axCbOdf4z97EOvjjMjBHT
+yfDkCjQdwwV6WuV+LOCvCPUt0y3Bm5I/TulxMXi/Vpz/CGGZPBsICik+qRdN48MuI/NG4RXZAbl
TC9Q32h4mrz81BpXtmABwyRrGiHBSLw1/lGYlcVEKtdEib95qiv37JdTWb0vexR75CCWJ7qseA5H
J/hEmW5gSNp1UI/yKfaD0rVMU2/8W8r2NLJuPRNwx+IZOxm3yInIUEHJheCaXRZaLBLCxlueLVK2
txE2SZ50vEkSYa/wmqiSsKN4Ro5nos3TkcAz6Rs+RfsKId9MiU7jjC8dWDy8fja/yGU/2XFRd7yL
CGBC/CtayvFqnvxe1PvSFkGwDb7v9ps/LPrj/8Bw4B8KB63saYGgOhFl/9pWFboCd5heDAYGpPBr
9NmUY8orpldlIZV0nb4T+OpSBLlBr7q/82qm2DKSY7MtmGhBHL+Xrwlye0RGM1JtrnLLRJvXbYmx
+RIR5vc5ZqOw8iXBye7fFBZ3j1bgH3fTP7900uw3vlkoq5O4b41HvKmlF7L5GstaFuaulUdnc+fI
ENq2SyDYmef38h0/d9XirqJnueqmghRTRa8piwHycfqV+acHT1+TYjxLhX7BH9iAonDyH3Z6Ks3t
K8VOL/EXZFQJ8LaXJ7kJjCbwzUmtNe3NLxP6oNdGE67oD+q+Xl56z3fnVa/AfMUDEAEC5t1DGhR6
VbXxlc5SP7bq51g121e34la/X5+UIWw7LS6Sef9fpcSorEGYZx3ZbPl6q6gYdS16e1CWMyz05Wpn
3AUAFhaHifkfyvEttbQPUC3zYf8mnY9TxCzcEBx/F57hQxoAtZMlOYvU4yocspJYwwhQh/E16sia
MWXF2l6ldAUuuGlKACHGBQGemqzn8cKapXcF3KH02oVfFHIiAasoZZbbZEGDnYbPA8hfmYcv6FmM
bllL3shWY1fRNa0ozKgibd+cw+5fWPlDCLFWxspUPvhK0bPO21AtRmwG6SFj3ymM8mKJQPv1f+6i
oniVMy/0o3qb/DTZvfyGUjQBBXltLvc4uv4uzVjd1SLojOkPT+UrKjvliIygH6QTW7td91TujKw9
Ue3Ehawmytjau/DWI3ujvv6DR7YzvV3EHofsBRMCry/GD9VX46gg8l0ku1or+N9S1WobJNUJq98d
rUv+SAlGQiS46V2zVt1tJn7v/vE5kUaqxNzgRa4ArL81zV2T63Z3jFCJq8F+kZ4GLliW7wlAXZHA
0P39v8+4yeiEs4avxEJXauDj1lBIOU9g1Ve+DL42Qbp0xuD04VKlOKQnOV93t+GE2650uxh1KkZI
ViS3knfhK/vEDoK1W5MeU3qBfVFsdqYAD83D0xiDC+vT5WC4UpKVkWi0OkHXjfPlxW+xb46TBL6n
6otVGNlBW43icPKFJ0GnfKo1DdvRzQF08doBteTnFnPYL4iDYalcCwhhvE3sJ3aR7cOObEX0mZLH
9Mcam9JGaFkd32zygpxRRyDArtJLPoYlxDP9jMy3FO+Yv49exGMwD0XLgz4LDZgYhh1cwam+WKBv
6qgmOXPqj7oSpE+An6W54gXhC9cdKHfWlq+sO1qTFTSu6+VTnKSA2th8fIqN/90fKy48I/B66kC/
2LFAQ7zm68knf7exHfOc0KqkmG2hwMLmkkhktPjvEHxoIdazbMRwLM6SpZCkNuISvfw2n5PLv403
3tEgoMqgN3h9QjmIl4VKwPeIUcJKZMOhL+384dxbCFlOtP9F0nS1YJpvK16WOZQz0c/33HOyv1V6
iobxDjQl6hBJXXxoavO9aNrjUpNrSMte4Am6EMdEsc/o1pLBB95VCSfFoRV+bYPDhGok/GhoOzSU
F+ft8Zl8ZDyCDRcpPLPqrAhoq0pRlcOomLRi+i6G7BSZlM6l3G0h1xidzIFmL4W39oSAdb+7jRx+
PvBWzM/FeBxPeur7XHWnIn+mVMrWve/hqZubOuToJdMa55UDc/yNDRJdNyhBMmxvX9Y8uuld37CF
p/VWFum5BFG6hfNPciwGUc4ZJBzOVJWnc1HkZkWiVMsJiuPAsCqqgPlDQNR/otg778HO1hP8ogwP
aKM6JCt55xlu1RzrKczM+BKgV3PKzmbrA7nYGVatfOJ8pSZM/ktx4LOeubQVIorM24GbcydBhO6D
dDDtVUo7CJsWTu3DJ47NhgA8wD/1RQqUvJa7tGMOR4F2QQL18Gbv7iDXobzZjH70dZrLPppu6v1I
ZN8UYZvhEDJWJYnUOH1FtmwgRWQhm2NfC+sOWu4j9Iah0AB9dpw7GACmo1k3biTZVmH2YWMw3tMv
btSHzLmbwAheycyGgC4iK+BK9U/0ZORd1EtDd1x3sd4Bi6nED76LzfIoo/8jITTP1aiHHzYHKEsj
lOsm5bQdUtZsdGgGa+MZR0kmmmLGPRQ2hIhkIXt1m7zWVyUtj9M6GTpOBlxE5U7mAMgHFkBEJMo2
uKlSoFN8wGQ6WOAa12wcGkOMmI9G68SlxB4WyWwlSb+IcxOnXQ5CQAJ1VPrQ+utSCm85/cFHZ+PJ
67bLsqFKga+cTZLSrUWIS8g32Zg7GE4j8erYcGg6uxJUnL4pXgZffiwiKBT7Z5yZvnbKpvVfRksO
4a/VosdmCy3jc9Yftx10LsKfX/9JBD4M8/TpMEN4oVqejBRvgGtUxPfkTMvQ/uWvpgMRZ2Bv4tOg
cpeCa8zU1xgcBes2eFy4tXqjLTYdb3hLKJifnvJcSIhLiAtFplhaualizTeIiXH/vCDgENrugXvo
5hudCtXxtJaPJ8DPh/uqCJOIbtJTvPVSrvR37tt8Kyeg9j9BeTMf15KSJAcrtWP50/pzFTDheG4G
oe1rqL5oliW5Icez8/RBjOMxTJdwIm+s096uUy5pdd8MMVB8OfwHhVXlrudDRaNs5/tJcbZxLe4k
dmz19Ji9QHXV/x3m2e8Umap3XAOXcebqJ19pR7cRYqsp2xB0+fSyikPRL0DgMFKek7TKWqkKaXr1
9uLedJRKuro+vqqpW/QEt4vM1vq7it8k1nTuNY6cr6KIJJJbcQovEUhLh4/3UccftSNOiHM6eat2
eZBNtdK1NHvqkteLHyQBYZyh2BY8xI/RwpHmm1sFHwO5ySMcwDHu4kDcjQX2mzI2b5X4BxeTnm7K
qTY/LXoS81RBW0s9UB4aYP3UyAdvjkcJlhY9ayOz66esv0L0ut/oDMcqnUQZO0Dl56EAsU3cGjil
QPYMQhmjLShdNPDYRgkR+osd2LbqosW806kSYRY/qlkeShy7I+76wIyLgwU5odJDc2M5t4D1qrzG
TRSADzeki19RnqXuDVNUTWMtGtOFZ68aAkmlrjcBQHJXuHqg9RrP1vvedMDvqVNu3Q4b9L+N3Ugp
VzPFHrYQLH3byYQt6Rl+grfi4R2AEk0JYCrUwzAn44ssqMDWWI/RidHT9SjUrs785Q9FZsFKWcew
1BHU4Af9aO+Rok/tGtbTPaKog+Eu0V+X6go8B7mJ37zlCd5kUXBLqCaS9WVGXPqN/pBZu/WaMcC4
6QgWYs9NOiwMJJjPKg/LOWF+tFjtgOsOGV4e5TJaSpkfXQ1HQMetZPOl5dHfHkcs1Fb9rGLggTBQ
wGKUfP1z+fyOiqpedd6Du0+mEY+EcYyCJxhY0KKDOzjG8YajYAib7HUReYxaEHsoWYni8a2osOxC
hVTZ6GeFutn1PN6/qneU9hJYPr6iMRPYN+xK4zHcjRvpik4WWSyO1/2lhGWJqLxiOihQWTqBLpwg
Qrs7GAjIQFAWQHOxzN7bCElz3Qj8GmEIMQTYpqsY1uwCo3+ABdS6oBcGFYK/Tk1Db5oT0BK2rhis
4CGn/0Pxzx03P6X7So5RUpagLDWtnR363GD1xPSk6uGIl4LFMy0VZj+zqzZ9kBMWU3avfHjjYL7f
JjuCSa7MgYNt+y/8O1qrid+RdeyrTcWqnowqZipGaWflzf9S04U2OVL0UjYJcmEVM2+/tGoJn0Pb
tBUJ4iygu3Q6DPxOD1F0AV/wy+keXw0dy6ihsixDIT0TorPIYAx4ObTrhZFnG/OFrdAVl7TxLxff
0mXRNWkEB4DJoSiHutYiIZwCNEeoi5kwiugj749tfUpjV8bCBcvIVO6Ls1i3h5nLAzxwMdlQnRbX
wdlE5Ctog8AwnpIeFtOyRTXY5NHt8pfJhwgp+YOb2PPAdroXGE/IF2TovYg3xp6whlK14o6HnZyQ
awuzOKpcDQDo8KfhxuiHm2lyLRThgIjArDdlzfWTySCCB63Ngw6iYidDJZblDEO13tlwmjyVcbr+
erAph8dimRJ0MKwEhWBgoQH+MvyXCjea56A2Xi6+EUcDiaTayO+8q5ZL+t9KYbDe6y8HmaJX4MRQ
DBXibcu503u+C1R9GNbsuhl+8uvSlKqUyQGbjPWrmXFZJuxthfnkMVx45nSiHR4T4QSnHGv9w5C2
baftwSDCH6hdBvIq9ZIFMdG21mu8ikFKBRg00sI2b02UPBddGk4OpsW56b2mhwFCtLGcNMsXrgO1
918f7ZVFgL6aeRwTMHpWYso2Jj/4bkmACWNLwbR0HkX9mENri3pyzGAeQCz9qlUC4r84/0TwywoT
i0QplTV+amS1ISjcWEAUf0r7b8+SYTaUY69cypPdQ/yTXbfYKgVYncwUyjJh20BwaREZocg1UBI/
UwIjRtStba4oQCwSklXYKDPYZxtp47zbkvLXKNm1DTIjOx4cZ7pZjhKHFi5ZFWLmoZLfoY0nKTkt
/q6/I3FpFpUjfkAISf6oohVS143XsNUK0MphbTbWy7n3nQPEUWHr+7tgPNh5feLffCiAF07QCmyl
LSJo+4Pte9uAWxMpOqutlXwNp+C1D+cwkBf9EIIIII5XMGa3wAKGm8r/yS6sZ0ofbuxXz5OS866O
SyHYaMHVwZSfbIftvaITV9x9cEkwc4ySNXSA6jttMfOSjYEZjnkxrnf9vB+8VMmmzb3WyjKmVsvd
xuijOb61uaX8nh1U37IjO3MuEQyzG0ys9uRTopAVbrxSOFRu3GSdYEzWLDe45QmyqwsuRYLX4vMt
vCE+8eEPa+RK+JKeU/mjmfPITSwkahQuORlTZXXX9TelLPZPX7L70OQTLDbTEZBrYFy+5GPCkndI
qkw6lOl+aVY1B1Ex3xlgWPM1vSNjqKekxEcV6oRyg2arz3JUApiufYeNwP/NR5ZnegS/9GvPansR
9+srpQjUjsg09OmqX4WiJeFupPJ8pI1kmFYATfqyPWfzfdOcf32z8aRRMDsu1UNloTgtlBofHEIX
XmowbGw3vYuC6Ev2jGyWvOPRL0t9nQF4TdHtrhbjYBCm602wQV79cXOA/znb4iJnHuMwnaXYb2zM
FOh2DCeb8TJ827KBaRXRIWVGzVifFvBXZ9KY0okJoomEeKPkc6PT3ub+WmUvT+0+I/F60XEjUWr3
HEqjcvmui0wDAOCgvLCLHFc3iPqONPw2gcZHRWh8FMpCUBwI+yYZejaE/l21h3O1PZ0F0EdKKQIO
RMvDhJBNPOxtyszxIm1nDExkMQQfQ1d9BnZMrLV4cVYwmymq2y82z/aLCnZa7YhhtWLrk0tyRu8o
F7RzxkT4BNxMfgBlolo43xyuu2lq3RTD07cV6peh1yOBmDjZ26YkGK2PR4TJg48orXm7h8bNBaVE
7DDMXw5bBAMSeyfpM1/AgFQ2597PVnPib/r13rUmSLRKFt4npvODSIhc4x9zHAT9tDH41q+ekpGa
NvABlAwBBnzY0tWCUhA9znJ8J6PJpHkEDEzlo3b3djQaOMrLvBXOmhoMje096rzPHJeaoUUXoemb
LOY8wyPV3fd5KXcJEVgvIS/4vo+5V9mlupGmMGqGs+PkALyOZZJtyTJLCMbfub5v6WBV7O9c2Wv1
dnwWbJYCVkfBJQSrHPM1slbHEiJpOWHBQYv3XhFHVhq66AIDl6R1Z+rhkJZ2WHbceET85PrmFpxP
41NaLWi6rmEal0wJO4pCQLjgId8S3gf+gp5fzJcEzunObsTUfaOBt9M3Cvr3aEg15Eu54xXVT8Pg
AWq6CQRwshD8PhfpFwBdSoVdWSraqZCwVk0eZqVwP7qjuSUuUwGRopOIWVSQd8aHArq4ZL6b9Vj7
6oAzLM+ylC3G1+xoaCCcq6QnuQlsurgizxQJmLoEnPGiqikHNdePunfunf0EGfAWiVo4vDzsCS0C
u4VBJpUWGJHrvlpIC9YDOcesqxemvwtd3memMPU99k1SM8+QZ23sYUJD7aUCvo+SKrElOutiwrWk
D8wUZb4l4reVWfqXFbDtPvLcmXV5nxn0vzXCIo50A+/flH4ZHH9WEbyVMas/PunCbbuV2yM6P9M8
BFRrkz0y33LYB1Khrleyfl5zlccswkc9A6ANVmSBreYJvawZleBiKNzTFw4bMufD+vHGyV3mHIDd
VbYN64+T/Ldz9l47RPm2NLkXaMQy+I4teeu8VnCFEa5mW2UWu2q6bQWFPFX60U+OsFD6/OUpDtyO
AOJMRqi7SnU2dcbIJKN88aDb68DkZO26LDjbzR+R7KggmAIzmpk9uyTNjAiYVv0oMkDf4ozS0REM
4RxRXOUSPc6aTLJ0B5X2twgMzMxHuMVLuCb8avbPMGXHEnAzDxKW7xu3KUaPHo/UQY6D3FQYyaaI
M4xsvndvDAIFxQ0mKBtmeCUFn5HR/m/nOKrueOQIAygV2mmu3MHbm/UvUAWrm9nvqGcPEzFe49+k
PyVwQkolStcnDQfnEr5j9tkGUigxAb5YrxJ+yZe51uRZJZkgGIwJSAR8DJCrDtpDxcWe8bB+tJNx
Q8tXYlau7vDm/fIul8jPHmSDCLPXOGu0SZJXORU7S8jLsz6pE7eipbsY49NI6rD9RBCx97FrsSxc
8QZ/6oMs9c3+/kmlR2ijzlvAomVuu/J4x45KH40wxfbESIguXEykHnNVqS+106kJs1JRrDOJXZev
YCmBwcctyAO8sShWq4TwF+hekKUfkO65nWW5GHYXOWPLaHd5KFq8yDQoc5zlgJL7Gezff7n5LzoE
TZ7k9CDFK0QHCDsOB//9DFUtds742uRmtw/MmDANua3LqoK8lg9Iq5xBCXZ0+GR4VpSH6Ar6UL67
RcKPtUSrrAlcOJ+E8DvnXXTT6eRgQfKRj0VbhOKyKdAnpB0DY7NpbxDX7wf0GugBGZH6Um9mTrwO
+nNLdusQs+4aAnDg8zhJg5ZOv+G2xUKIUN2amSlhJhqxEJfpFS94kSp54L3zMrVU0PBQhV9Teqnw
SXziq8TyCj4Cwfq0l+l9zQKeHtqtGudWtKSrbx8TA/D16YOV5rRhFDz7XUSHs7UhB/pK6UNEaHhM
LJQCq2RiaHoo4/ljLbxMPS0Un4O6Wqtx4/ExLYHjzTFViQr69/A20tURhqKipxXnzk6Vn6mFUtgS
OPxk66s+wo3IMwbzXVIroKHiuiVDixysXV/GA1J42jZTlY7oI+WVgxQkwc6AYvmQ9iDlTSVpPS8t
L3LjY8yfP+dI7qbshPAnNQoDcN0wRxoLzQXQJ8ppMD2EfbSjlaaP+dOlDqCdXohYNwEcyB0jQjMg
HjqCanMMhMKLA1CVdu1eRaXChGIHd/1NVmxc2d129Wj3WRZERiqo0GvoqexkQe/x2SxNuqwUUkaa
WVGKnpnIooSIHlnWc0ZNneyW8peOolkFm+S+i2jzS8qCQmV9VuZFCpfQxELwHtxycIyyqQnmcQVX
T+oGED5CKY63XxrGqRlafhBYIZbuypeyc3Ijqmr7jsk6U8hT/yRRZJKXqmGVucYBN85ztIEFueql
ANcR/RRrVT826VHHmOssMAfeKxMOfWRYYpH1Tx5gqrXkysLqG90KYl5iI6JLyFw4h7dmGpjuK/nL
OB1UWD1lxCi0r5eC+iSWC8lTkw/YhNB+CbmDedXMGKxSt4LsiTbd2r+0eSU8QPqdtN6n8Sg/W93H
hKByx95AvlHPsxV5eY8mwERV3P3PTxiX4v5mH0zt0we7FT7EHcRQq4B1vqSq5C6JvbnvcTJaGOOZ
7JBIUqnpD5pdnVH64jerWFVX/NI4yGoDOmrUalN5YgG02e9ZfO4qWd/lvx0hakhwCskUxGQmZ2ja
2K3XJalbzH4AzI46oP1JF69qsOhCFoBP7PmgYlXCHXrosVnyQLtXfMFoUOchmlUTpsX11lVulorL
DPauAv1VTNRqdexePE7OTMq7v/iIwu+mk8+dJc1HGIls4PP+b8dSC1sys823VFrURbbGbEj9z0tE
kuCtNRCBQ8skRTro+sFhIEQ4Y/2L6HtltD5f9ZCRSyRuFAmzPf2EnEddIdDzk7zHbczDflDYKdZj
oUAn8LB4VahypFfc6Zy8IxayG9n7Z5AZUyq5v50EdUGdzhJQQLpY8xBTwU9g+pIKC83CO7vIY03L
2DNHVV5XktLxxS9UbCTA1bhZbFOHxN3aiWogAvBcqs3ilQkNUjtuClTlLQ7uVxY5m6JFBfIv0Nm6
fiMAksW6ly1F+2ZWwjxHhWGgdavaXGFlauoCW2VUiIQ9h3YOt4sMHC+SohwrLw0D2jKUw72bMqVj
+Ye7GnJ8MgOleMFAfsrIUoSt2LMQrO/oOnJmGFl4ThoSwopz1Y4ZxVoru2R1PNuLAYDbEPZd7PUy
OMVmXDiQjmKVdb0cflSSbxbjyUgvTpBpWbzHh7zIfV+rS/Qge6Z7fskdQGNUGSCsVbVPtvinf/w9
1NKQF/QwPPgFLM6yWlcxF0abCz3UyfrXtpeQy/ms4y3gKC7s9Y4X5rRlUeV9vUppDGnqG9FamQIj
8LGEtV5hn+0zX3ThTNcH+xAlsZvQir6R+sPrw6jookbAyD4JOk4LolXYsEcu4cMce8/hjeamODpp
0T6ZSqFCd6SgbMpl2Ng6X05x78APtOcqhfWMhcPmFAN/0X0DCowgTARZMxdg5+ndP0mVU8xXljYT
E+XEAIX875M9o3nByKnc8/NrodQ9jmVdc6nHt2X6ov9yY6bxNFv98Nl0h4kD69jex5MEJc/QYSSO
688+Ym5mCYIqIwj4SS7foKsWtDq/Nx2bUKPdwCms65udzZCfrurgRCnJitzw8QBRqTJ9h6SQrsx9
/HQaog7eGyn3UR5F7PP/yFnHiVr09d1INu9dE2uoY3b9rdU2ldrWGOYd3oZ32I9GtM5uW9JpNZ7a
a0o0P/YUHpCVYNPV+AXtauSrnxkQAQqzXN7e4OdlTyHLmaAPiGOGcnLBAHT0tHd+2/fnG3MgLGq3
JFABYAThTQHQCuCuT5peWIcn5YAAtwWBHVenedVgjYAAJ73iHav07QK//moaqesNyGNP2aZfT2JC
pnEOHI87EYOfla5gBZ/yZTdI8y0B3dBd43XCZ+kBRiNPL1b5t5pKhumccqARAzZgVJ7kdjljrDUv
hN2VAXbgA66N24Su18+RMfGC/sEy+gqW5erf3zmSSlniSf+EjapG0OrOmdPej4oLce8KsnYS8iSa
nv1a1rgX4oqh79eymMMhUWVh4Wo59ZLrKhPK92nQ9iNt6aWWJijyrfjjCVjwWAg1sN/ZgeQ8cA0a
+pxVqPWtbQII9yx3RWrT86r3if8J/QejlzpXrDT00r/J9TPRsMyJI34dRkugNRMI8mc1EVs7yrwY
zp1IR4HuvM0LZN/uF6HH+gPPDaIeXgavsENt0JIv6LWXtpkA1oOJthKawltKD9HzaoBl7SFA6q/K
rUIpqawt5jA6LWyqHO2Rhu9iZqbnYHVVoN/8jSOnyh5xyYT+PfyrX/qRVAaMGmh3e54oRUT0iArG
uMlr9jLBqHIm2bFGpR2Ux5WqyoyiaiGEIFuyyiWXg30oowMMCsq6f1UpQTM/OcrLjTMfD2kthqxf
khAOGTR22zEPj/hx2GwppMj/iGVc5Y88BXZ5uXunApK99yNMt+jBiJNzq8F5QLF9ULKQAVaOF3fQ
b+kHlKnM9d8CSC3pBVFmtCeML5OhnkICvrxyBRpiG1Yto92ubm4k267taIV0SPpPpkp0eXg62ATt
bnoN9NT5jo37ki9Ykhb1Wcy8eQz6RbCUXcrr9YUdifdj7+laHC8hU3nMuAdGi96Fp4PuGu75IW2Z
MuEprOSb2NzpfCi3yRxKq9UIeq5LQTBf5kjCvjpXWIG+rsXlbxTmZRgI+4gBUs+Xm//2v8C/Ij/A
fdp0VU9TpQJQIpJ+JiDctVmsmrR1c5S5vrUOL3IBrb2cYSDepqMJ1CEMfSplTRqbfwYSq2xFJ8xO
J5OWOKYp4loC2TVCq/Me4oiEX9ZQhBGZGOy3hKyWK0vvzdZNXkZqEX+sHEG44sHiYsL9xfb/6zut
u78r4O2OfTZTDMsrPTZ1MJQh+bIWeBzSTndp6xZIpX0HeNVhpQ6vGAd2efYsWEs8YZYRsPHH3bPM
HPNAvbkGYIyHNYbwe14gTZ+MqvxDfXI1XEo6g82XZMhEzU0MUMFSN4z78ZcLvrGJGw0haYHmKwRU
0Dxwv1VL12oct8TWTty6tyBp8TKbYUzVrIUfcidJXOqeab9MDMwG7rwu2NeyCPsy9Jts2AWxG0gF
1xVZQPGTMa5PQATw+86rlLHpkFQt76dol5AcN8o4LJNSc3EVmZ6x3IIRIiwg/VgC6KRpJo6yy2DQ
bWGfR1WzySl6r1jaTnH/zhq8dmaet3q1DSV7+4lfeYudPkuUG3WBOmvm5RSPON1lcRqsYvEeQmiq
iAGX2wGkQtb4zflUTmm//0Cx+prcFlWeFEXoALyCvFbRUfEoAjklsNm6v5s+44tGlROqWa5W7UcI
lHw1YIuyUp5IIE9nEG2cqycoZ5gfqMSGs+bjNraYsJuUoapkkZXHqmTdhivA+rqG/CIcYEizjMTN
CUz6YzSgR37r5Yj+h46zXw94nbqh3kSkCcxS5El2Y+aP2qZdlV8oIc5E5JWFquHcqVnGh+/2XQ9b
lK2TD2cX/767NNMyiMohgxCNXKC/6Pcb4OafT/AbWuoo4x0/gV/7jz3SR+3QoWhP25Kn805guZY0
CRUuq70WjBCfbkuLKZfbcA8YgZ6XAa8iwMpTYHQBxX3xuJk6QRlFd9ogPpgUQE39ZnAUEhYVVgS7
jBHXlY4VmkdbRxBZF6pUMTD5FXIVVn5mb9MxM8Q9Om+YrV1o7nwkzzcE6LRWgXmmTdpjoF11CdsW
3+06IjiYuD0eecQcoCbMY3KWKnCWDrOfvbM3Il4IS44OcSFnhZ6zths2PxXMoZW8pE+7JNTy0eTR
WXWm0b2q75Q5/g7CWbOWxPnkFbQFpjyqvTQ0s+5cBfQT0hE6aN/uqEDlhFs2U7chGOhYAiGndboD
wuFyEmVCPV9orWRtG+iQAPeCTZsLcbknOKdiBcRewwPb2j2Ey5Tqp5PoRKBAdwU2D0zO7qCPKM9+
3Nia79+xI3SogjXpxJo7kCSaYPkqM3+JfXtIY9wCOfIRrZd4nOy07EIE1GZWeaj+hcYciUUpkyS3
GxHytDuCENqHiNqMSh1MO/IRvzBMVaS8ECQa91m0HQrwlISjV5apVRCl6dHpi63eI+9hTlOGS3E/
fzKwErCrOPcAKEXDEFxAq7B0zickhyDe8DhtapxIx6xUe5w9234pAckZ11+W2oweAn6lHiPn6an7
5/4849fu3VjbY+laI54nUmf2TkxynEAyCPYjihFippcozHiUpAbIMjZbVqWugzuA/M+t68IOZb3H
Y7u8rvHYDj48gMEH/fglJ6U397cwwbMNezGnzhzGTCPQcRZ2uZ4u9fSc7/Kho+o8Mm8osexhmZAT
/ACxJ3ReqMn78DmuAXAuKVHytNDGQZ0MKTKrFOcAH4EbyOY3Tr5ibf8v3PgAyYt1tn5m5MZ6s1Fd
4X25c5+hyVHKZM723HWpNMm/yMJSmTOWRb/EmoGHik9/aaAEaisztg3mTOw+oRt+hHGB8tEbHpKd
pCWg+zLl+cG19j2UIb3708O+x2JNRp2PJ+x8RDnH34Cj4zyVl89uT2eCofESHbMszBVr9ZcX6kms
EvHLIcxNbJvvkq/gMk/EyAa8ZGRzAKFke35z0TfHUkwW93Yu2UI9gu/0VNm7JR7eVS48sInEi3xc
2Dxb1wq1ctcxWt8wFONoFn30mKECuG53nCMwLgqTXQZVCcePUBCA615opajwyPs/sMjCfKz3HX3L
0zn5dCS757Un+eVBmyAq/t8qcoiD/AD2c2oDUy5rOyLpm8UoAwW3Rvh/PlJGJzMo0i0OJp0MK3UQ
fHGxHifrrCVLlPwhFgTiSDqpHot+KdR5p0rFagarCESU4Ex1zlyJrSCbcilmbyO0CosWeyWG+Z7n
YlbGpSbfqsKE3qsmgdcozWb9GOZlG09R2lTc43bNjMLAghHn/qWRGyvz+iQcbRkH63k1LCIRVnXm
ScISYYS5ziA2KGkXe4CWQXGKjKcLAXUrWQ/S/maocWGO4xRUe+t8kE1DzVP5/RqNM2SqHUMoP+Dn
f8PL4dmJnTc0zQkW0hQCBkEgbBVxz11ensyzCFv03gcfnngVa/6DN0fXa8qk6SZjbKH/bXcIDfo8
MaE6zaF4HCvu31+wi3SG0Lf8OJHkhlCy8wNY10yUYFxEu9WEB2qph0smKcvuAfnzRrGYkd+UvGVb
ZByDx/NthCfsjIqvamxwWWNaQg0VIifdXW7sVFNu7j2bCL/fBVo+gi2yIt9+bSg78ELJeMpu4fJ2
IAbHDf2xOkxQe5k0+bY7W1JSnS0pozHcZs0qknRiOtpQI11SSHXqQHbkuH1et2Bk5p6OLWAODnIx
CEIIOG1GqnlcRuTykop31WAyhNTsb+u7YVh9qR/0NXSffCMQMqGyPhApI1uUHig1JDfSGzvsOuYF
eN6sDDOFnHsuA/GePlYYbLSuXfOcpYFvRwK/bLLLl36wHnaXR8apmG82oHDGHN0cNWYfaVXeACvo
hg6BbVtqudo1sas9XrQ93CVE3YBZsomtPRb2nQusZbg5aG6IvNws0hmuyWwuLf9rX17B7LACHstY
KJLxnBiRC1CJnObUl2/xdbqjMgq7cBsU0Ohzjr4NrO38gRiBZBy7SDBgMXbE4iUU6ZuSNXOQwZ0b
QYjnSH5bv7kM4r9VuNE7LYDwN/VrL8+kf7Z3wjPkxL9gVIEoIM1PLb9PkobdN1+n2qfP/7c2nw4m
Rziym025hzDJzOuTgVjKX4cQ46oxcaXWQmh/IQNjTtXBvMozah5yKsy5SRgnMtf6YEKkrQz0YAQq
QXU3fZcuuZt9uCKuK46Q98pG5uUAkc43ajtmhCNwpmQ/hFXZdM9Lr6FFYegtd7WOYf4A7Knvmpc0
fWjatHeBnkGU6MphU42hAp+PYJKlPq6DRYpTUuJSRnNTmYBzhf8dSTHdfaPIKy5APza/rgjQBHc5
G8sd960/HZUyk3JzKeS83AdPNQpj6Oxszw2Ih/LKYKsGeWN1slTeuFY3/01LYNUOLw0hoKFwJBfz
cpc4pVD+cVggypjaehHrfbXUtmkED8eqlr4APYtd1cvtmAcQc++fA6LZPLzAuGk+YHuZvzSXwS+e
gV8s6pCDnniUZRd2xMFHo3YxFxii0McFlmRC9tkHcW98XiigATl+TBMoFughunW9TdtM0JKuNklm
4Nqh6SfcA46tHru70yYbWNdr6zyZTNwoEwmX+HQdHHUCrmt8tPEmF5L+CJM6xxN9XT2yYUjGpnkb
fFBpCH+OCeS7bDDRKopFH0IU2UaV6wTYx7rhzLMEi7RnfPQqfz3lSLUa55Z325p6hCiUoAVF1asd
7jcHJpuYfoE3SaaCihKSUvJki1tBTf/xMc39WIJpKavxUQCGvIrQRswoF74MBLppZUgZeRRLpVf0
/tR2/rR+tc53aQWvhe7DeB95b6n7Mc2zOYyxbJ4OLLSBOUYOPH/uORGAGr15DbqriVdzzdaz3/io
Os/WlODYWKejk0wZlNpYuqnnWOdi1OwpTGiOGl3JADoq99xaFxdRd1OhHmWDPqEzYsjpa8pw84+V
B04NVgDjOmR68v9vKkKMlq9e7garmj/ZPMcOZs8bSgn4bTcthmg7zBkrvZwzXo4lKpz+W3u2mcZE
URF9tgnwddGcjawc/7k6eyfEo3fc0/Zx3FBFilZA9GgUsf9xLxN//9oh1F4k0mLDoCBVu3CdAHd+
kYd3zb9mw+T/e2vNAN+lvhmNvvyLjEVyhzCnFrbrsWS+ticy+T40isdIj4VVoDkzFhAXUTMTB1kt
rK+/56VE7C3oNprCO9XthpJ8Q4wOTQ7qSuWPM405Wa1aTXB9OrkC30WYYQwLElL4U0pqyO1Xwhaq
zzquGU6eydgz/vWxkLtRBbQzBKrDApqlfKSxxSJ8FMKvdMRpTmLNdo+43h7UQ6xbzaEjt5rJJ0hk
e0bhZ7Mo4nxN7KxhLlwfHRJp84zQV8JdoUBfPQNXtin+zAAeMLIO64JlwFFC720Lu2twXlyqnCPj
4aMplUkjxekIeJeKWkTe987bQ1Rx6Si10BeY2hqPI8DcmlXiVZbhmKnydcBZrHggDeDbtfwt7q0f
9ZznDvgXyO7CNTeb0624ZPeIfCwsXjS1shFh2YT2Z7jmGJDF/swfaeyanNxSs9nngtoJnIcZhqVB
ijf/z70SUR1TX2v24lMsrI45lmjyscjoB4gOkwvvdGAmx+d32Snuu97YPW0zi70mslo8RGbuukW2
4LDrW4bX02D9RWJGGayI97gDZkdNPXFQo9eOSCHhkuxycI92ylbCHQ/exAnRhGirI4x8YEwx6/vC
iXNwo9sQ9V6cei3bQb7kj4OrD9VzeoL+5AXFD3Teo3tK2map1Ry6NpOYP5YdrnqEFBYycftaVQ/O
kH+cyChQcA7/N2GIzU8s4zPFvlOXkaHwCjQk4iMBcR/R2HBeYjB3mN+QRtl/KYSLlJc0I3RJuay7
4S+Mp4gm1on7SbZxiPcwrv2+u2CEr02MQYgBgrMoCijniGqWRCRMCntIlGSYSwxkzaoYDToLx4os
YWQquoHJ5AlyqC7olkOz5Q610QEAZvhJ6NNqJuab9+ROtKPcN9bMQo2WCoCiJQbLgzhjA3IIMdc6
KDYJJTfEn0WE88IHoHHGkvogxsURngtcaApOhOhYALGmZ5Mc+vZntK4tKTa3OzvBlDD+o5wty97k
bIIWM2pIJ89Fa8xVTtR0+PNKzq56xMqDUtX8vyCUJabUegIQDm1tz+6MEkUc6d5Et8ruFBXdivc9
/wplR25TAtqDryBnsd6bom8XcxjmjUuS4enUCN+FmKUQ72SO47om6FThM50lvxVUEUSs/qqaSO5w
YrOjYKx7h4UfGPbrI6T/ZJ6brFOuujcwb+YFk5SafTojCFiq2erI21eQ+vfSAG+jCb4h/UM+fmQZ
YFl+/lyXYF67Kjr5virV4kUcJTE/x5BkM235f94huublsk7zbTJs5njJY1UAct102iQd1CTAVRRR
V/QTJpX0ZhquUZ65UVL7NP0em89nCIrd75+FX1LvyYPBUaLslYAxJ4v4ydduqgw/qAoOT5vcNRUI
NMRDeSdOIkvgHkA142D0MZqO+Ms68UO9ZtaBcm+4FC+obCDbgdQcrUzidE3tFC9b9eDJyJzcOAgt
u4a2Yb4M8PnrGZRLck9aeCoRTu0rH6911hwld9FKXGUsq5J5FAFwaeaqTQBIy2pzWF1e50di7oXd
HUwlyfp8ALAVDmrZb0+D8LC0xKUdspBrjMFNKLPhxkbCQ72s8Z9WGxgyoLsw2+fCUMGKjyW2UoJc
Xx8pLLDtt4EYtg3YzD53Wod55QyzSQZrwGeiTWytL0eR6IIwJoVes0UDEkQUuLfnVUUJgdOFGFLi
0J5oQfzJ/NiJ8VwcAEiNohCWA9Wy6p2mglKk0E2A43XDqmECz0I6jSyQDAfD7jR1NV9Wml9B++l3
gZcpv139SbxXmcU8u8TVPTsg/goTc/7zxgoeiFmGLbVwto1Ed54CGIQOfW/LcZspfjhb3LG5XY0q
RR6wFrt1KeTtdcAgPxWAfpf4GWtDB1A7q6wo9EmRpWBypY/vdTELKvxLvP84en5sfDO0sd9R//c/
XHt08hGyaNWa3lwlKip9dqn9YH5ZYnkoYxVeEcSR2ybrt7GTAflezJEQ28H7CEAgo61uMlI5zMWT
EeTIjmhyHaGOE1kGtGWw0wI5BA81J5rlRQU1irU7s2Iq3NOgUnVr8N6zlTzS4bOs5k7dp8slkPOc
3Z7UzYggYi4HKQqmoAyYmaLPslfxR8rZ4/1y+9v0gMUiDDYtH8xbxLrroG1qQKqcKpWrBlOZVAUN
6FvTZva2y/CUnL42NXkTMdvp7M9HlFzaE4lU2eidXrIaSz9Het6/VVEHnpbY+BLv5RYxQlfEHIja
SDRmB3VhN3b84AcOBvGNP58atfCK/JDQKtqnhc21MaTpPcwBwDehuLEb2l5C6y6DQ2uwsno8faLH
QV0ebXOglbYpm1ijNCZvFSaltKc0JCB+tZBo5RhvJ3FM6j9yv6FnBXz5FcnhPP1xzB7b7OG+qi5s
wt0kTSuKspxkaMkg1aTRb3jvAnNH0x10yfhIVWwPsDJeFSxZOFe7wM710zBwoleotBL4t9lh2VeT
Yb8Mzhtc4DfQqbyFvVHHOKwjW1M2hIe+Bb9s98s/5Vq6hQ2LW0Qf2a1LEv6LYk0/ZbWGFPz9yTvS
rHMkwnYY0z/3S3OKpFECrO3K5uBxFWHER1ZM8nK65lF5JeaBcD9vmbm9xAG13pkXnz0ZJ45rBCUe
Srsgm8HTwcZHXvq6aZ8W+HQvj968O4OAEySbh5k1CADehHUxF02upoI3iU88vNJykTyos2/uIakj
HpsdAeAnHs40PeGXReRB4Nz/vx/RI6GhKzloD/n4AGIF1vkLONoPQFeGVcPhuvONEpy4q1TycDPb
CJ30crF7AVRulEijvvXZrODKv6jDtrxDaVxYiHuzh1iBSXDlgLOJ+b9s/6JYozXux19yuDT7qGCL
xrO9M8URPcJqgM9tdoNfyZwP6dGzrCXfIbait8GmMY/w8gsmMAwq8wvgWv95vHdZXFQEIDbm+KRa
p8HDUyYqKRKWpfl0R+GECnlNsgvAD25UEeeb45aEVLqILI72Z2/KwR4OMXsTeJbno8hZROJpPO0c
3mAV1n/W0m+5PnTjlBlTNn2I0K/OFVH/o/19VyDdXrCI9NiX+ksc7lRIod1EnWxpNj4lXKBCqICA
XKGm65Fn5bebUDN9OEFg1Gfc5lgj5aq+ES/VF8uVwIQzRULjf7mH+mG1UqXH6p6klUI8QEf6CPnc
j33hDjLeZjUaZyPPc0yZF2edJjxBSckuH3xF/HpyYoXF66fN9FGAKQQTxtRNAYCE3OILwGRXFGhO
X6gZa0G49Jm01mLjTLxdRZhlb6fEHmqNMD5lThch8u5MwXgpUfhZQjQERsnJvdgbzL/YnEDkWY3G
gb16f2f+v0fPBelRrfeMdEKyPy2tGDjfyy1Cfb4QhbTYIFbsaUz2jCOWzzA2v4NdF2dcqiQSUKSj
SRmwh2F1Fr8Gqr7v9C3/bBmz7sI+0PUvoYqDay5g7v6/HRtUji45gFpYuRfMSTT+XHwUR8qts8FB
XLYOjtQOa8Yj2wc4C6BI64GTt0opAekYOXP/ezrFPgX72Q1EKvXU/WMGY8PkC5BR4n7SwCIGBLxZ
Jv9LN6IIpWzksEfDCdBiCZ4vKE972ODCF/P3yooTe5zY6ZPeku1MuH9rihC3qNb3LSXfOLJQu2YD
6ekOeFFjuNzX4O+c7T9rbdugmgXqZ43q+5hf9eVELNBvAnQqXV8VabkKlch4dI1UUbKu0U9P8F6H
8vVaToQpriFTAnL8z9VJdYoDJZExWD8xattSxj4+lsQUHk+Lp/bMtagGmuWIK8d34QVfrHpd+/UX
pjyBKt652tUzeNblF+MWnZw20ldICmAzoQ5Qhc+SCEgdkYWQMefXTpuOgbYWA94zhzg4n35j984x
jqkIjVwkq9FFMhDIHnb/LW+s4EF5iIpfybDwI1NzbWEbygoffuLtmTagPoTnUusUveZks4c1GeVc
zkiJsOckybim3w+zOs8lraotIt0g5odXxxk+WIbmU9CjT346hTyzPNjeukMwmfN4NfkXolXptmW6
I+3ZPFlqktuWZFl5zrSBqxwgNXXC6o/nn08FBNxM4UQYnBv7ouWSsJUQERaAiRwBXGJgCBmf3hZ2
q1UboWadKmVDzFmaaTleWfGwuKywCxLevA9ZzfYlTZDA2DJHmXu1Vb6NcscU/MPEjljXOsaHMQJW
t9xgABiWn1d9yfDgN3HkPYwsF6LoSMWkaBppGk/wnXp72Bs55/QkCuD/WX4qpEfEBYzffIAMimXJ
nMPFOYWwCLrJo3xaX/7UMH3hcgV9fX8nAY/a/nVAtRZBgSSUpo0pwzQJ1wsltv23Ni7fAGbzAwfb
p7SiRl4pzLMFb8UepVEUB8JUnrx6qLSBX/4u9DMm52EgU5uaGDoORDkj8jIfxg1aAEk4YTt8uzQi
TOeyxthF7CqqHje/mMokjlz/92dn2BrQ0GB7oEfB06Tmt1aFhYdUKgTzMzKIIEHO7+s5xXkLRaSR
53L7azNsVxmoihm9NWog4kdip8bbIh4YSLGs+bCwB6CgkTB90W2MzW+9bQ2dLy1OJVkhprpTeV4Y
APzMK5tdMb2t4xIYBjKwWZt0kThkuYpntxNI0bjtQArceFbZ+RoaMqfKEadF3vbp4zL3rbg7pmXP
PUP3ZzYS7FLixtKlilhcWCHCgnIfYOlqIMZhm47mx9rTTuoAKjt/0f/NeJd5ZuHRJsDID6goMFtE
9uTeMH5c5BTRHrT2gDByW7iZ8zxZBCV1ZUvJfhQGrJDVTnUs1XELGRTDoTSvmcq8NndEmNX3THHn
CpkWDmoQu0CAdxDrOjkdc6H6KM4/yJuGdnXg89KVoQU3uvVjlhL3clBIxln0QdEErdIek+QGHv1F
wOZtccYNviAAZOa1AC2f4NI07jhK6JtgdRPg5xgBSTNxM1cO9jYEzTUJ1TZJFHL2gkpjm/N7kuaY
8XXeT137lfS9x6ayLNFIgV8AvW7B8+ZYI8j0Qs5sRxnmxKD9ObYB6I2PSZNOFQnATR37SI4ysL4l
dze54x/QZYhqCz2CvfLCrHnmP4RXUM+unnCE+aVvOV2qlhpUPfhyZlljAwmVKU2l3uOlcAg+gJ2J
8rrqkCIsdlbQf+LAeD/SpC+Y+ljwVeg4j/e2VEE0kViuSp4nTpZ7JTT0BQGJMBPlB/HAPWCOLN8u
UubY3krMk9jZqGSzq3XhaENS3CTAMxv6ldsCQqXDkTzFSnVcpskViY4XpXjHj+Gaw/fNjWRNohBk
5afVTAtb3oSwphoQlaXSMcR4IMVy0UvU8Z73dhuxEToKceKE1Nr0mSFzOxmyHLYWJfp5xJUILGxo
y6NJsKr8RqBKyJtBfiUC5yn5g9Je28puos3nqakWwIVIBxRSx8TB3DEPvegLWeT/Lohq3Pk+93tG
z82NFiWIStT8RktT1gRcvu8g1UE1B2H0de/Wh+i+42SdJC0YdBsmTeEUuld9nxFF/iuLoxt0BcjV
Ie/OWQO73ku/OtqbZbxnl+J7warjOOmjZ5UpXl54WKWJDhhmf3SlXRdkaId2ogsUPOrVXAAUD1zD
aPT9yGToniaYV4DDQjjcGqiu5gZQnKzPlHiejf9t3knzhZTzokrvzSWygpYt4mvTuZEEV5p017VN
U485ouC0xrrxjcRabiPDaFTP70W+Ov4TSYuI54X6hf0c99yWUmFUHgttIjETC78Sr9U5lMNGVjbH
CAKZT+ayGl+pX7CqMnrpKo0rooDrm5BcLOBy9dpIg/Meo7gmaHBSKhU1eEpBBOGzsog6FOWVey/m
p0yAhrgM0tXGTVMKCswvz+GLp/Sx+oB3j73xodCiCnc3BuCyrgXhdgD+PsAPlhHNm8RdaBjBF4Gv
eSDLomxudk3BgvY8JkiUF/OS0dj7wuw4CPeZV/cN2ixh1JUv11MehFBReaby7qWyqbkFwyuD/dBf
fDHplnTvJ9b4j0anMHSb9i6EpQe3PTJ5PpjfZhDWGXkExrxbGPq9iNr8IJ7fKXKF7Ry1ptIfw8T7
Foww+ClriLcx88GmZSHBHs0c7luRpYVBlRZidkQSEemQv43tz0ZF1ZvVZVXuFQCcxyFMutp3bzbt
fnh9M2M8dpRXcUDe+wrsx8QHJQhakWJgxqwJxao7Ws6Nk/2ksiXipvFfkJeZtB2avqK4xZzVyvpq
V8sE/CmnofmojOfDAjGKyLCL+7Hd7eXX2mrjmtyEGDsgMV6kUkfuUcR3QLcWdO9+pJ9lRwNw/9Bf
XqgxkMEM12LNkC94maeenaq2OzIoBImJ9xNN30ta7VAJHs2vHgjf2/PFPnMguF9OsCUjeOzQ3/LQ
r/AI85B7IVvfGDyTezUi7Yi081tVhwXYJy1HT2vhSVZAm9j+Q2Tt1bsZ1w+i7ycQHpj7PgyTQ8S2
apaVFaRPxoW8g5pd7Omkv+wEZ2Tfdv/peY76xTZdRRqwesbnOvhDkQqSrCbqdScpUvUcnru+B4rT
cU4DGbO9cYxIn+/IHFo1PwCSGlHDW6bhlUwXM7p10zPBE9+7U38bQj6yI0VrpNUv5Z3UT4H2qOIc
52lbP0fQ8/rANXiht2/sOi1XoiM1MRbQ5PtpAYOgsdkpKxIuskEv4zJJgBDzaX8MEIVyXrTEKcmB
whCpR7vOO7uI7xgRZIdl6fF/ZmJZiGV65oD+g+8+RlL1WOyMad5TFcT4ZhFMcyXn07O7FluTENRj
lu5hfB2CPz/udd5oUz4tAxwd5cyQuZx1wSGp6/swyOTLH53Yq0yPUF9jbbzemegziPHo44pzjQhy
arnz049R0UrQyK/MTocbaTYNwkVb8AzsBuD8wa9+tBl8b+yVemZbQNtaFSqc8Jri9N10ZsZHtivb
8LTAoLp59xYoWfA349bNe0CGYlg9mZa6fjYoFebjj80V2LHFozN1UKA6QV6v3bcNzamrbXLQi4Mj
6di2Ss0V88aAo/EKZRF08Suhk9TF5puDqU+v0snV/C9fVYidkBkXH1FzRWrjSAkZGgAZPkLpBFk3
i3DIbx5YE57u0gG6IZAGwKv2WQaoKIja0jrrxZsVy8VOdru92W0lafraFkvjd/M6m+YNVKrbYC2x
oYhEQvciGFWQImjeVq+5MIf4k44C9JbkhndN4Zv6SwxHYCGIcn73thTL/nrcWUFCvOi09uDtBlFQ
ldJh/Kc7okM29Z7jdd0pZMj33I0U7bVe3B8Wb6FsCn0Oj0U4LUk7JOXNZD2orMx0HVkaCuV6BLs3
xmHxni0kEnPgVvlTYJdEkH2P/ivaZIJ9yio8WjdR9Luqrwq7fmwxn06pnwWy3p3pmjZGytDQhO1E
NlBBlkB0YA+13ojYjB3ibLlC1CAd7g+ASuS6zECvYgq6u9KTiEwm7NCLVfGxcHLQyaD2BtMOen3f
AWVjsmMO7op6YviV9anCIrJnGBT1PQRtxtD2Y/k8QFz2J2LVsPVI/xGXhlV5BsAWNqdzE0t1sdtl
+4kJJwp8aM/DDN4f361vh2DbPngtjvljshi+ZSDlAZIQq89PmIYupostCP0ToyvXFe23520E5lC4
DIxyzhW5ennhAoNEPuETuRbZ8mm861PBnBTMZKU4e1nrgOg/nIGRvLWjX69A5BVOQdEH1WSDrvcM
CW6NJKP1P8zqH4zewF5Cg1G9nHcd9y+N6WA+WZXXKlrjLXD6ekspemGQfsU3lnW9KuT+cm/tzCnq
xwXM7MgXonVWcedJpW82L1YzABjfSJlniwpb5gEXRZVvak+EVQEucYa7q7i6jIasMEGR78OWd+z5
P5yYQjDDRtKfveBQ6jMuIfy92F6q6By5ilF7cBEg2vrOFdnMdrDG+WD6EUqt+5tpg9nD9rSFFkaZ
pktNZP4zdXFDt+D7WSuL+2o+XXzOSLbZfVP2ctr0tBRCDZIXpkwnedbhu838nQwxS+gLaFxTuqul
edsb1Uvr0516+EiWXGMhes13FToZWQDw121EeGe1GwgrH6jrODixI8HqnQSU0+AcrkTMlpU3V59U
V+KD++C+J6xELLynYJZkevfB7A0T1H6zitSLrMakXKSR+eR8cpuAWDC5Ye16mknXQ/ni/KGfnjDe
GCTbSfkKNT8rvQTlDHDo4l8SNDP4RVvjGkirTn18tO2vstrgXRxODN7eixfEgJTHbfVFkXDyD16r
k6BhKL0dWIUVaSwATAHN55XkdzUF912NH55qoUy5KEhkx+dGxMSin9RBYT/sO5TduEjajG42NiOu
NqlU7YAzJtnOzq8opRUKf+nNCkSLWhx0HJQ6ehdT/MkKNtnToFkb0S5sCieONDlRMTdbXeXI3M7D
ORRq3w3Btrfvq4Xn9HpcTH2nSZ5k7NIfYE6DUn64aZtKrESONgTZ+ez/ijL8yesWxnSoXjYfKlF2
BpH2fuWbFZdhZdYMjebBHQDMn9Ei9DlwgZI/T12tQ2vBWLxjL2uYDumq103gt0aH7cEeZ1x0BAd9
DLEvstSLGD4vSirwe5uztsTH2WPtaPdyP9G15ctuifgwwEmdlyuyPl9g7gw8RfiBYLZsOso7FGVs
FINQhDBUyBfm0xY1bCw8Xz+o9chcB0unxNL+iK1Ci9QnAJzF0oO7vWggT+vX6TOTiMbDPzNwMsRO
6/YNuRJ5yGoem30KVXxVwT+H09tUxBq3aqL3nxFaEoKCJoyZFcNkbvGnsCEFR1cS/RNprC5zv0br
R5Iz9GmXqDX/JzIJ3tAsIar3gYUzfDWLi1lrhDw5cn/iSio/HtiIqkdFKBqLDBGKKatQ3009k+cF
IGYSfny+2tShQf4zKpq4Ai8W7UTdifO1vj79QN103ZWgZyotz2g1Wor/riHwzY6sdrdZaOD/Kh0T
7mw4BmUpmbE3PLYCvU7Rdl92re8PC26voHAMSmwMoAFJ4PIFmn6vwTke8P2wahyZgWY2ZPqFrvkk
qoYdgEF9MCe9cuSLMZ12LdKImKxI26Vc1x6n+HPc14SAKbXXnmyxqTKjyejgYSJWSBYqXayP35d+
vvisJcp6lOTjVM6MPgwvEcyGtZYz3iAvu0oQWZN9CQ31AzT+Vcow94X6EAtNBOMYFos5bAdIzjfX
22OVCQKgnlnNZYNnwAcdMLWm09CS47YDM/ZVutI6sPHw5ucSexkkms3DD2bIqdlZdIscPxkb6Jud
IrY5nt8Rf0rOXn0Gh1OOn28AKUX5WDtPMpnCeqeHrBJntp7dSkOWPDhV7xItBIBw8jYOYufOKwGe
dlJXDLh1BFcYAAF1z3QgrE4jcOGOOa2J04AmjX9ZBHHr2JTkjECcyWFRnbeTxW6FKT4OA71VKVtK
ozsxsR+HWeXM5UMtS5RGhmVp8Xrq6U3PspbPC67W9NjcRZC/JWmC6BFj9Mt7dFxcYnE8QY9dwIP/
eynVK78flEkCih9R/+ZawdmmH/W6WzjxBpq6CR2UsIxnqjxLPnGVAG1xaJyUeUlDYp5Cf1QtrZSu
Y1KKuMvw8QfEfcEF/oyNxq2B64cpJ6SP/PWNTq5sDbFENiR4aR7B+KkZTbup+XfU1x1e4+hHU3z1
jAK2c9uji2aw8DI1R9PMZvcK0Zl00Q6UN3g9EiYeWkWF/TNYQX4QUQavYmulEfpVvbc+0uGv8DfH
nLGyMM9IVdePzWqzaZ4eabH4HddWvfEkJM+SAdWU4YsOoUh3cvCc8MjQhmE+P88fynKP5eS/uEI9
Lvnik1NeAaEa/Wb8O2C1ASe7QLv8FPxDFFNucSVnZtQ+QN2D60EHfNJaVsPlv8CUFcZX1SHXivLu
ikF7F0cJQTcNWAFF2QdigZAgayQ1wysoXM/oJdIORi9WVXNA1g5c409uiBiHfcaDSKirW3mSr4Kq
OClUNYETaYU4n03vhuMBs9AaN3xPPhmMoZre/JjQpht2MuSVJ3gr5W7mZA1CgB50a0ol19dyR5n5
GL7qC3bPT7pbfdmSOREbNqjGmHsbute8GorTWT+NfPmWEr4xiGBETqpcDUMq7b2l+PF66XTQAJ6r
bKXycPvfp767M8QAr2KXpnkjxlLbXECk1yJT1TSgwsRnfEspFJ9uZLhtPrxEknWS41xQxOqB2i8v
y/cuxOfVEjoW+RY585yLWxz0WlYvkXWndxQBQjKpJhMNEhBAXa2M1Ca70pOzEEa33lmIzRdC9BqA
Y+m4/hxgflwddY4ejiGLippXywDlEzUhlG7R1hgvvg29YDN3CoXdXKDOTbrreZIRrQAKQgXu6V1H
D+3aDxalfIDq94KQEeh/BrhwozenvgHS1pAVkeGBhVyHU8Bvjo//5BaiqRwfXil7iXIRKg+mhBOJ
EAZm58/3IybRG9OIVXNwu2HGqyMQgtSx3vtejer881FY9qiTSS/1CTedJCpWIf+7pm0MjvlLtHxy
/5KJx+p53b0jts5vzYHJ3E8CFAaoBLH8FfhaGUT1JEH5k662ov3q2PO4o8smq90PSQTB2oVzYEjc
9NzWg1TIynR613cyRkvRVZF0YMczzzm842duMPA8AFhMcKBSPCQiyzZz3PkfOy/4r7cp+nCGiI0V
znf2lm008XW5knfgMfl7HnRQTdgFdUwPLe6FWV8nk6yuWTTSSpuKQ03XIMvZ9354ydcAB2n76KzP
UHBbappycf1H07o1nXKCFKo/g5oxZOLzKpfOy5rq9F7ORVJw/e4vLD4075QZCtAB9PjVddfbL5PT
x0xfQyAAMehA8yOCSRB2JiCu1S8k/F0zsJuIK7n7fC5O3M8PRySeR59g7g1MGOxMMUhqe8cPoUHz
TPN7CvZXkAnDUcG3DmeKIzdMjyD/k2dqdh0Zk7twgv361pML3hv5uuJgP6bISkldQtSE3OBZ671S
txV4CRk1YYU+dYfmkH5ovYIykxw6hWch7lAdNa49qzlDCyxr6gRdYMLBrYcgV4Wb8oF5abuevR1r
YJzkJugaxtAZ09f5Fn6Suvy4huIbFCjPwYii9Ui+zYmxlxxOv55ovyTXamCI2kOV2Y3xSbwMVGi1
yWFB6dXNsl/CIAdrx3CRlRWxa1UeLtCrMIVGqW7qfoJbb2Q3ye80apUTICzcVFN19xp/0wsRjerk
NsF1FpvQJo3XhTKKaQS5UNM2VCkqg0EyL9cghD89HowliZ1k3Ze11VfzFqeFxMj0zyRt9aQYkAf2
VGfbpyh633y3gJUF4blcNXw1QaCqI/ivoyLA+jXfLEOdJ/QT0HSEbxSywQjB6hvS7H8G7LYhaz69
LIur3gAkVxP5e9lh8084kLHq2BrjgOgq6s+JwqNGA6KET0Mgtz2DaLI/y1EM9pSe6NdaSjufGjnC
qs1i5e7UwWgiYTV/jODImYQmkglbamBTlt+WzRZKk1XQBoVKwn0PGRUlMqOw8Evsw5wJi317qRlh
49DSYfFZYTewowGme7LdkNKgMbqQSBZ8ZH03TnPcOYCMLgHiKXV90Vo4C9YV0N2ce0KqVvovENc9
XgidImjluePMBvGpudPE3+hk+PR3e5j+Ct62Kt7gPboiLFL1dTau2v41W8GchbkGE5Ki0vTzqgl1
vkp9QmMQpY2KNNDxiWBbc1VgFkQSbkRggNGp2SGlnSRks9FN5eEPyiVKkiNYbLK1Aw0RmgZJK+LI
364vC65Dfvm4gOfAe8m5p+cDCJLy80e/YWLhp4NmNjIL+/9YMa9ybZvT/T0pXZlg26wdIvAkDDw3
OfEx1NlPh9XoFrtTO15BNWsagwGB+zbPg7/gXrYjjD3au4urpo5TClXKrZGlbHBrZ/10qdvIwQ5Z
TYc+tl21iUec+Hv2MEKtsPVPHEH63SHelYb26w1qXM+aYqc/AyDofc10OvTq3tZURatapia4QkFD
6XFE7R7iDiq2M9t6O9LSWGUhzlx+yAHepQMPJn+IZX22rIFrxxNSI+3Ih+7IM9LKM3/6hli1ca52
cflEXe4oQXa7omFMG/z+Z1bQwn2f2ocG2a3KH09CeMJfzUeSqN4vkbHY7IoFCW7/og44rx4BhXpY
fjlXvn9p4U3Qu8mYGMTgg6DK8vpXeD/3Ihcf1AtyIk5YPcbQ0r97oP4ubM9X2f82Gn1Va0YMS1DC
BtQbMqEV60VGpaMu31C0OPXO+t+vOsAvYcu/EuAhBsz2E4sUuTh2kn7K2jj5QAs1S3WwzwVlCVzQ
nRuMfhkql3wsKxkBNIKt3jbpabSQwFyEO1GYe22etT3WhNNuNbo/zUMUsXOTVnaubCqgoyQLXUFP
59RDjeukk/Jkn2JH3QDcXn0QSm1GhMFqBIxzxPms3HzWvzMjWHgYuLB9Ses+TGmRauNg/UaQPirJ
LkyFCmJn+l04Rl+gl33GYCeHI4+n/FJ2FcBm+X8E9iuSdxeIlgZdtEI798FzVmY2W+objQrgKjVT
rY3U5cFdCWmdzUISxmfqN8+9BGrGn9J5v3yFTETEHyXByACQnTAZyJdYRFkSiqONBGuj6CkNGH5v
VN/RbdsTySRiL3TeksfA5s20eKm9w45XYsnrV/8PlK0TEitxq3kQAZpP7a/T+AfOxGmoEJn2B1EF
2PTz5am3bJ81Af6FMyYNKTY2uqixcVAgTgxg5MlBNyI/BLcFtPHabFMsmlYpEgiegiNtOJ3vDrhB
Qrsnd/5Qfr27S3VvBrS2nuq9RI5Zbi66IXtZ4WjPmeehidP2BhIG+X5HdyTmbX/+ntURw9RXxDBO
0n+Q8Tl6xXe/8xDWglgR8NUSW8R4IAyoFHRSBhrOkmpcWC4azWnl4PotGxybroBhgHUMHFu5U8cJ
KTq67Z/afbGUbZxZgwp1QqQmthbRZi4zW4EpmgK/RAWHhw6FCmmPEf6nfEPBH5zRxRtA1MQQCtrg
ysEmDi+ySo19rSZhKGu41bWuRMl59viQid0hzbTbRxpstUBQaJF7i4rGeCZFAmkNo1tgftIjSh2O
wSOnWci5cCmsonFkgiYiUOi0Cw1WTmc8zUb5l2S1lxSXAZzQwZR069SBX+TGOVVK0Xpdlx8AF8+e
L5l3dZwxm86sHIJlvMrDXU/V7eJVp0MYIgzjA30E9UtzPWIDtFeO0DtwqMMk28uDiyYwJLTzOC4y
Duulo2J5i/w+V2TE0TBwt+ZFpBbf5GSvCHEnuIDxId2M5bV7gVrFe4Z/u8atBJclumndDeHVbwJS
CcBZD+Cwwvv0bqwOnEhpVdRKzIKwd8IsyePItiNDnIQa+vIJhCyB27KqFAitGhMfTH+H1gXRpoAx
uma9lCoUVCwQ1RNaD1KcApiPGQxbpjdN9jTrdRklLvsVRhxV86UQGr6wTQFbGmkskLFHYv/Auxzo
m5SMaCCfUXOSQqQfp/ssek1EEwARc7Nql1d31St3Vqv/WUXEU2ROQa6lkbJvGns+eaXDkaN1Fy0n
AXeQLanQYmkEN3Ehsszymuh1RcNi9OgsV5InLPANZUXWa+dDaMRiqH/2d/S0KIZRC+zMYNR8agNT
64xGsHUV9YrrhBIansmqYtIu3gYadJzR2xhfnDwOYhqA2OYvQcoC413paNYpRAohOTEvgznGcgA0
dxwz0TziOLTIHmh2/NG08NKAdrgYgTNKv3Kag/SCTFGcapN9dUhp9rKzumyUw1eGMxAwOIjcTRtk
Y6RdF8NSb19R6vNa9992ZrwkJNlu4Da7n4jL1CjBgwqCXX0iU84zoOD+sO/DhMWUz46Tbmx+7LTD
W5U8O2xZnap+uQEcIVWVS+ddiAf7JZUki/I3XDG9iqjWfYdoJIAzkaBrpXRiFHYN52zi4UoAYQNY
wsUy6q7rgCvts9pX71eEk46Gbc1ktmD/0XbTbN6iEbjKM0YJaFoTfX3l41atYbYQAxHh3XhJyeUC
nV10rYpZTz5gBD/GVEKO5P9cZKqxQjON8sJYkaoiBAoCpVftoB6v/vsQR4ri4r7k4G9GgIkalUbJ
Hm8gWB6xnFipSHGS3g96WgpIPvsgb3mTHECspcVcUwUfPBN47eWZrfdaYXLJZd4Ya2jSJyg/py05
uHCvIySYUpb3C6EevgwIKG0+7DAH9lWAnty//+uGSdjemvGSpTtYSX6otOo/RUqyZB+t/QexKiHv
7xGD6Ek8fyXo1e1ZgwCh7JjPL/hcGdOe3teyI/VHbCaKQfTTVNqDmM4VqOFzGvfy92sYjZlNhlkF
fr/tcVBDmOVN5t3adZS8qKz0mRHZR+v6gk/KJghqcj/4Nw0l9be3cn3NLBxoI4LFsq6nMzNbufHF
mJz5JiORxo0gpkn+e0EHQuY7at6YGD6gnQiCUmXyiXQB50HI2mT2zrtatzJpp8va4EEoWHEeFYFy
89FLWnxim//E1cY/biNXv8XH0aVNcap+9b7Agq6JuPLC743jE/R4eprLUf66m3mW/o5Fi/N5x6nU
wc4NS/lc38fy16YKVSbHHMNcRe30GmyoDfNOyWdNiQXiWYR5cS1nZ8xilh/uf+VYtQITVt6Gz7VZ
sBiIXvoSmpNG9IB8tvcbs3JgnR+yb1QtJ7EpgLpLv5FXzBgKR8O5TVDyMfSZ9L4p6dt0tv914Qle
ul7/+MZ9BY3v7tKM/7eaPk5VZb7HzlX3BPTyBRkgDh0hg4T0IGbsUrMvRsk5UPRy5j51d+1CNC98
v5eVlwtH6hg9NNam00v+4+RTKdZpvfIy1ZnYl3D00oxNWRqO6RIELaYTikCNhv4tlS00yFKzC7C5
ChFScNnXfU4zDGBjXl6z/iLgDkE5qo5FoMWWjPZYqzvVIXLhSbExNIwfFGfyZbI5GIvNreULX3zf
+6/jVS9mgu7CPZMquCVuyFbh20hSrCOVhgyOZLBfnOVrsML6Ub++8mYGAgB8EHGiAaP2V8VXafBM
IfbzuwT7c7028A2ZEfAvcUR5tHBu9FIXimyeBLH5Py8oOTZ7GoRVtk4WPjOJ3SX5TDe57PlH2MER
KvkxvdF5uyFEMwkYpd8ytj2ymtRxVJIlxbt5yqFxjdsm6TUfOMV638FJpsUjhMV6z6yx2rjYKx1G
zeALuPI7Jd51XA8+AprKyZ2Wpu6B+1s6mGdeGHMKYleeaIFn3CPNm5RB8x1e00xcwjQ4r4ML9Jbn
Q29lTsDMEXAY+rtmKA0/Z1atNDJIlBl6OscpGJzRLKVVlzoefKV8rJV1RRGuXESFq+/zTNcyI/nd
lbu5TntSQHxDD70DJ0yu+5LIqJuuaLVtSAMiZn4xYV7xzSoSXqzhRMZYNFWJD5FMGA8NmIolTSTS
CLvrwQxSgyEfEWzvMTnqpVZ6PZyuIhpUodSGjHwNz/eaWJK41P74EUvuy9Uw/650KvA+k1h2kE34
NFNXRzEuwbcY8z6JuxXIvnbc9SfC0N/GHz502PiHYcEePQTZcqbazFMN+uXdgELsYN1hjjDC4CB9
9gjQm7QyDkRYBoDj6oM+YWuLTOYq9l2ESDXuRV6kTQQ3bkoRCaOxXC/cxOcizEeTdRJIgO/tqEjm
c3jTm12Skf/JUR29VaA56RRWcEIPfLhs9SRy6nkHsT9HLth4DztnEgJMiRWZyST7xFaQ83BjqouA
7qkDTKgHRoL4fMCEoJ4TwwVWvDB5l4sZmCesIq+QJA7SWIO0Q7txUGSWtEMLWvmzCtQxb6KrEpOE
Jn6roaFqMl9vTT+3Q/FwYaJZ8anEQpw/i+ZO0N0Qh9cSh0UpLeH3kYxkB0Pr/eQ/kIsukL2o4KSW
Dbr/drIZk8yYlAGVOxUHEbraNhlNzdU4eKyfkRceFA+uOqSIaGI3sSV6Z0ud7/4I5cx8yXjXLs2P
VOU9bU9OiEGkf8QFaHYdpvSWQN1OHVfSOShl8o5f4bm1RvR3jOFUSjJSY3PtHqbrQa3wW8TyI9zo
8askEb1mXe5B7cRqkjxfGLZZJrWTYB4ivfpR5WS/rpmTQBGO/x/2XfiAFEu3z1BR23WZ6cOBBYUH
l+7pMP8P9b/KDdcq4G1kvZ2mCoYRKKO6VwSmTsFjWIy1azbjHOQSR4SKJXefsXvfP/03mTCZlAZF
06vs9nlYh40avJ+3EyvPTedMZuNVMqUMYmshSbt9rdpebSJWoMMoP7icOxO95dqrb7dyC69db+lv
kcPYcb40Ge7JTM9g+PkOs+4aawsUNSJpWEJ8CC0ooyMJt6rupF7ZolMdFJh5ABH5VLLziILkJ8bO
ViprbTt7F87Vgc6gVfLjWGqNaw0QKvYHQC1Uz2+kaQQxx440q/jPWAKqijSKlNYaEyuj4e1v79v9
Ol159ta8sD9tfjiUiLPTy/MMHyKd9wWJvyhB4YLuUZhoM7DNBaVBxEFZ24l6CQVsWHzZbbQ0zs3A
sbT0hXeA4zWQmPFD13R+nPafBVarI828oQoLfG00CROpUEJGdbK7os4166aAFc6qf0/dngY2M0Wg
3wl+RQxD5r+kiCo3T+YqaYe8QqpDwNylxoBF5qVzaXMQC7+IjP+MqnCp2RY9kZZkE3zXIiGWyJdY
EwpMJd6J/fDMmZA3xrU6Teq8+KXWq9ApXYk0nvvMwcdsFXPGt1gw7ucLrnp6OzeXkYcQPT+Tc8ai
IZD65VE20KKeYGGEWdkDPAE0vW7VmtpPeQy6W9K6cRoEeL7ltzFSOjEAwvtb7L/6xTFQSkrB/AVt
/rUNLGjuapU9Cdd2XRhc/QKlyAOaAkavKssAjLLc8XTi4yw4euECWu12BQI7xVT0vOQKQox9wj5F
g+xtJpVBNK200R3fA/37o4nTDK1AZfFKFKAip30Yfmgt6GYar1J1waLyY5JTweeGh/InhClIw+jq
vRqW2q1C9MIpD+S2/k6IRA+5eim4e6aWBnHSTiJVaGZEXfGmP7WnfRqBZmoJzvCJLk38Q4dSh4Gw
mkyUbpQq+Gc82yRyM1t26CSspJ8osYLHerclVTivGZrXF60Pad4KAhCdpmoxX3TqADGd4S/KynR6
Dys0uZ/88Tmj4uJJ/YdBhML9t5PHfv6vbxEGHWzxVUrhCx1SzoJlv21Qbi6nrNCXpqGJaYQDfsI8
8kRwMLyLlp5ZoC7azqEtcyN9Baq81hi4+iUMMYZ2bkCRSLEZsaSaP2VQxl+yKh+GJNGkuCVC0zOB
wGP2NIIvYaHXGWBdTGJEXHXOS9Cyi5NWGTjhudKxPevxMTrfPNNfCWNGadD+Gw25HCjpT7Rdr142
4rM7uxi9ueIsy5v/tuMrKG2COFdsiMpLL20UPmrt1IdYdadyVnehkjnHyx4sgjZq/QTLsd0XXbVN
Kjy0UmMAoeGxRU+xfi8UAnVD/23FNc3cKfGPsbOO/O9NsI5KhaejMcDsDBCerFYjMd3gzOofUmHU
/2YrRBpY55GHhGiEMhgho48uAvfjKQusZwX3W8cdu2UedmqGb3DMx718a88b5LxsLgdQTJ7KX/Ix
Bs6FEFtnsECErWXmTozpiTzt989w8c9dfpnuTljMZrp6Yon3LV6Ea59/aN/gUcmEHwqBMqrLmkqo
HtLDU0u7PyevMBn1Tzg7NNbTv8tGwo079Y2wZ4NXstdQmCeCZvww9VdcXKbkhG4UM4aWMzXRx/iT
729+rsLvZqKPrFieny4+A7HsbV7d8I1tLHw3IGDfNQ2UVksVi9q1+0tjYOlRAUhU4akPXzrc+YwU
O4zyM+5i4WkD0UILmAR1ggFr1BS1xHVpsHToLUStIrpgi1x4bAcShfB51psgrQTSc1MVBndm6Yc1
ygUNctVNMY+16nd5X6Vk5lNeIIJCS+Vn8VabRb9UMpdlI4LoE3cqxJyxd8pajWuS7Pxr5GDb1wc9
5PA6uwJbfZqbAsudkJYUyq1eg5RtuLZObqeNoff6bFvlM/yDimcDuiFdHdRNQJRxtlRESTLSjFKm
WZ+05tKKdWzEBv+OYlkLYZsYgbJ6VGB4DjdUCS7MkCqYe23kTVqMOSvV/ndg71UAanoda7XeQx9w
Ia6BEKZnBRhK4pSrlBFhJZTHdyG8nLNOqtHh0mRBUsrEBi2OP2Tti1VN8CLDDrfrz4qhKwtrfxDc
1D704EatlVSIMM8EFkK1LJwtvuE8pXt3XQIdV+KeQQYIOCdc7k5tBbrcDgQvVfZVc3ejuetwdK78
rSNx8AXc6CmOi2NZ9NY5QxpjUXAch5f1DWD01G0j/OEZlky29MLo4qls2PTYwrRQdjv1h2JynGJs
A6p2+7V8HQe8YCF1QV4q0MfHYWBGX/o5wQSedTE6fQ/eVpSrMWVYwSw6HfgA85WOq4v/SuHRFTZ1
dN8d4SuH3M8jaBXvIYiyFVuTwXxSc7FE2aKsmvcyAl4iXJ7cTrBCifqBPjmNOmgY/xyyqbol5FXe
CzPfemcJyhUZD7CTyejzJMWUb0C08PMCowpna8aLXEgZPAeNoZecp1SW860cb/wYPuuCOYnW/L/1
AZXdtXYuhyzMoRAE7nBP1Wq6Kf9Qe1q0rENuiDHjwVrt3nbRJqD7QkcdDy7cjjkPFgxi/Ss1nm6q
JCSbf6pKF7c+kVvBNVbH/7btWMsku4IWy/g44TBPsXK5zQEM40BWLwHF7/Ag4nTSAe+C7h6Gb3qd
ptA8a5f9IvqBNRTyMosF+Qpq6sxPIwfeM3kTdxV2wbR8yZij+6hc6/oSbh4J751vY3hhZqc86Cqa
OZNIiXGgUAD8Ge1mKcWmu7/VeNBL1SzBSricBgtXTLv9aV3GkpWukThpU5AR2/mLTDSY2Ojllpry
UvrlvocUaPDU+Wk/PWxa4YVisaWrxqB+R4txYmkEMFLcZVOW8uFA972acBptdIJydnIlLjmwCaZD
+HXCHXIe5g5IvS99mFrwF2dFUhFeHc3yxs4ZRRh3Pd3WgRYwpb3aYhahXopZlD96Lbuc0PO8RSA5
0Y5vA5AZYxL4Qi9NYmEG0VZSEcNVTxg2Itv4azBwICy71h5E18cXCC6feND7V1/+CnVb6IhRL343
FezMlFLH6E4efl8UfsRjgC9l+ndYTI1JBN5Z74bttrRgURRoXiRHedOhsSJ7/zxWgdbcLaDOwApA
0gV+awycswQZVbWhmUDWQnC30xj6irFOV/Omgwc7xBho12T92Rhw8lZ8sS3RTn+BxdgnuSBEcwTt
fWG7h7P1F9jq8UvmPTHYTEmsKOWHz67vbK8t4/Avc23vaPO1wRPKChGhnmXtU0a8d/nJmgHmsEzG
IQlWZlKO9DmOLye3n3vr2EsQw7uVylS3k9LLpdGKKbQY9TS5cX3q4rViDURNkRr3R49hZOg1u9M4
0ZT5GdlY+DVwnAakhdf35wafiU2lDKf0mMbkDMS7t9OV0vDpNLhWufkG8Nnfu5Idzws+OARy0mJL
wiE/4GSMV0AA5LBD9/0HTlkZGXPboIS77EPbLx7bDv7ofFjuT2bOCqW3okcY2k9GFszp/w0hYzCT
c2rkYvamHuV64vvqsvRHqBjrdexRbOOXAeuP3Kdgd3hBvy1JLLtdVoRVFy05ws9q2vENlsPKyopm
rdppBy1IqFoqF22C0myjadFmeNxxLLuJiG9hXXcoNVgi04+KHYtWosLL4Rk9syqMEeIhIwbFiyG1
DIIGwq1GKzI+4ASkEoC+6+9SXiuP+3Ho5/DJ+2qUUda+w2vQ26jV33ZjoYnwhBNePFKr7QHuW+El
W7FoceC8JWYg87YcXC2G9FhmA9X6xZ5PnPnRawaxbdmiM6w9pZA5QzgTmcNLPG6z/sgLMTQmRNfN
wbgBJdPmnb7fZtVxiAJZSWbN74/MQVEZTI/usU7Uun1/UIKmeCytl2SBxQXeLZ4Fms0Y/6cg46d+
MDzNOKm+/Kkto8zWPQ41WGlbGMk4gGw1Lx8HddaXHDigeinJQhX6RLIXlVgiLr6PC2g0lBGf56O1
jHC61ka2bIPHgEa87gsDaZ6aKHtTdNH2oAJ7YBIDgGuLR0AGPyoXDeVLPVCxkt38IQWstZcB3f8/
6otKpMSXiUGypU3fVJFUMqtsXB8aR3j1IGK1Ho3HJV41Ka+yfS/FjRaUAFgK2MMzuiKN/rPci8k0
hDrvlW8pFL0zmoMkTOYqc83Py7T/245M9UXgekrTHkAYegoafbnLQSFUe3yIilOiYRcHWGYGxOdV
x2/ftTHx82OQMs1UalJFq/W5wOBTUX8cx5JxaMQp4Ro0l1E0Lj7FijY7H/Fanv2eT8OCemGnN8En
5MMBfuxJZnKD7B8Cmjb6izT6ytpMdUIeXg0tV49Sy5vyGtw0eKKnome6JdIciVS/a0NS9rqYVYeb
3KdFsjrsLKwwpjhXiNScFEIA048bhoTQ91VMIta2Zw9vw185IlHTI6XBYFJUfex/laSWN7AfwdQ1
6ifqQT49gQqJidduuRb925VXf7Z+FiUPV9YsR+pXevyXO7zfRQCCuddunEzQnoWH+Rde/NZ+5Kos
C3cNa35BBE1VtZdgqpl0S7LABFRAQFCYosZwUjcoArZXBRRjVJxQ9q7TCIn5/miNt0tDgk7PQIFR
KZawMTJOw86D54d4I7o0FbubM1Y6LffNdJCG/H1KRf65vbhvv6s5x+y3lzO0Hb+AWyQgrPLVYuJi
Sg6JNTLQ/9J+KKrXsBm0RSZdOMCSAsb7Tm4C73b53xbl7mEYnC2YA0GgNyW3FOUsKy3iYOo4BXoi
WNiH/9wpSzSDHreBWrfTHNi54+U13EcDXZjbPaanqpugPPW/28jqFWQH1Fx1o9jAtGMd7JwPfncp
OmvzuoYBGGiOoSPmZWrlzo8rtv9aOOTjwanJ+F02ADmZGykT3/NdXKdaGsUHb9WTaiqP2rXqctO3
3vGAhiiCs0+Pzz04+rKxqsyrj4vloMspSV4Fx1dQLBAfRBbEWs8sgd5E4LlCKychcRFjhj6RoBCu
VA0Feo720b7w1TZ1o0ftZSkBj58vXa/bX7i6PdlwIjJE6AAinqBKl5wzbJhVrXugO4Qn8gDYwlXy
74/D6RGbjsMiuXRVHL56DrlsiBVVyC77tSutUNB8lgvUe7TKyDyFflp399e57uQVYsRWrW5gQClj
GaIa9Ga08WM5uxCQEVt4VdLvcqEuKeytigUR6FuRNyvUSHfKslUaTJAWDXfnzF+XYTFZsll/qjK6
Ue0h6+2l/x2+tIl2WMsZ+KgNdInro//dr8NIy9Ac8vEU7VVMQPZKf2nO8M8AclUXI6yTwjHBuM5g
WODGjxJFUR+BHI8fhGZnRWGaWnCd4jbGepZkwmGWuYL8f2ruS+1KJDRJWvJ1DEI6fgkhiZ0l8FzL
qWWea3H3sTMUNdI1HVwOM0iOFdoVwy+PWyd0v+X9WkxGaZRnIZ3ymtLsB5aGYwpIje9cdiRzZa+J
ZAXbvhLEeYiRN0Fj7QAT37UCJVrQYtXGyjZJXLqK6tBmsIWYhu0cNF5x+FZ63Mg8M5vYGPwQ/lG9
MID+0lOj2sbkcbQQCNS8jNH5BrSvgzLAX4eUaU/xonxTQTXg6Kwni0/jaead911iLo2bcngZPHNv
uhcj7lyjJfO4Q9czxEqDrbP5WexmtqD5daOuuVa+J1B99nSHFpf+db+uCvSHz3YUq+QqT6q4xoOZ
+uJAyLO51stDL9FtoEtCZlL25qOI/KRj6TZpwIM60hDWlCGY+pz4mFV4n1gGiXGLREpxibbcAqIH
NKc4k7M5NhQ2NcVWhOT1c+fS83rUjajdY6hO/cykX6rbKlwDFOdghUOJGGsyG7pEauaguBYBr0Zi
bIlkb+cIS19usOa2qffNAL143X0hCHCrivrbdzcd+VRnP45VPefgJiHgLGktFhABjL6QVyG5+sRr
yhufWBFIW3mBLCrlD44+geXFYWE/hiSddIein2UpVF+1afxfvvRgkamVQRuTaXqM35VvUDF5U4xm
KQ1g/EIReBx99U0dnEo8dPuhZtxEI/bfYmxDwjdPzZ6TKqS5i5GNxRay6HDYtm+XvdLdkfgK1P8o
I9AAN4TAShtvi2zAzFYxC0Ns6qBbd1QKHKzlquEtJx1afgjtDiN59f0YwAIJdhMwEf14owiOKeOd
Zarwn4KSfebpy6OCougGtHMgSC8alN9P7QG1ms/q5pneLsE2mY1jd0oCGoUpBqukMUl5HGUszuHt
omkzFOlGEpLkHqajYIILj1l9VTclfs5O3drZUudH6udg0AOFBa4PnOJLHaU+JLmk2xBqmsws6RTE
m1FKeEtMK2rhZQ5ZJ8joXG0u7aZGvhVs/vMFpRcr7m06AhiGnvXrnfomuyxJAuV0iWa0yZCn0d6b
LEyFNeh4xONn8noRKgeGoowejOQabrTgLeC7fvEXd3YUkeTZFeSmNxm15ajOcpTFENm4MDWBNgLm
tPsA1DbDkeBji0E4LOpszU9rEhU2vQqw9HYdA43IFOiwZOh5izc1bMRuhDoZxo/JcXXi8v4GIHjZ
uUmr1l6jFhdtPn6U5K3drGsWTczhYRuOD/gDRZGeSgXX6olt1lqpW1E4ebBIjTTU+rSZ2Ay6pOB+
jik8a6fqhdy0D68xPXYI11rBd9m9XlreSC6FbPQKzrXR4bUED3WWfoKUDjwoA/jpxcN2Qdh4wnp/
3og8IDlIfxm94Tzuj5V2A89Cxwwk6vefjeXcVF+R2HZj7DAE9adKk8S1UBhtvfWu0DkaqvDgfNbL
T9Q+qxmA/UW2tcdNDwa2mdtmIZYGXlCxnKyRzZ7MlIPplU5QUXuzRQkEbSCkzhQTyzs0Q/tGpkIA
3KUVNbUlknRNbgTD9mfWPN5niZ5iRW6x3Pix17smgmgyXlnDmV9U97DSSExTENIEPiV7zYBeF8uR
O19qqryidP33Xe2GbSpmpl7f9npws2BCl+Eq9FVKySM1dGAFYq6lBY7te9Sp6LkXzasalkzM1bw/
HVL1LhqpZZqVq4NXjvizPRdRg8XBny83z3CQYCmLsKlIkQW8MnK7O+1CwUWvv4D/xbju9iomSYUe
pKxRQDG7F+aNoltNhBBuzChptBpQjI0GMT0fbUgVKkecomRFcZzfSyoJCXo+vgMud+32gwYZy8MV
kmGt9Qp6W+tolywMAkeQ4UzWlZneejCFUz7xFdEv8HgoBSHKJeIb55r+MIJL7xLGptsWfJLhcWVg
QqeYgsBBoYQYVNgIquw2y4tl42bUTvhgWG9Z3oEOom91rsNrcG9UOVPk8PXA3QIjcBYUD1cNkjDG
vlwAPc8ltsywBnfUYEVWfCdFRQO09MfZUlvcFvT36Ij4Ce9TeWDNsXBKZD7rxURAGMwxRn0XiX4u
P9MrbywYTi8rMNaEDifxZQIHbFIbWq6FAp88uTGgQjMWBo+/kIbOIibCexG1ciM8iCvAbmTHODFP
d1RV0zQbd+dANYV+6LFRCSYwl8A+7q+JVFNHZw8VbLgsn30FRQ2e1Xod7VhoALHkSCwfIENUzNbq
Dce3SZL+gUD52wSeMAbuQTlbSC0tpxp/kRAH7dSBP5uFIvvSGx/JTmwKUZaZYhVlAtJZwrhdq1jh
o4gm1Cd6A2930/NTd4sx/Hes+ZcnIgTSnsdQEgi9fEO8ixhJVSvxvqeBxW+p9kUwiR96EUPseBrT
Bhi3amp388cwvAy261fhRTOKb6fqIYNHIx3i9JB7rGhkEHpLobIkh80N0YsHFYEBs8luC16pH5pe
qh+TIKxe3O/Pi/W0SvCpst7IXZFz1nDEIkYAzRUr0J/bQYEjYkAUM6fFcbZZ1BIWe5SJYbhGSNr9
FEyazrQhNGhOO9BUd2MKCTTyplUfBWkpGmhtjSNFsLgz4mP1ARO4OVNTEQBZsxAivm7d8zG/ygu8
wKJGo6qeEGkwyj6mDYemScT1FBeBOl0YiShsF5z1UY/xzNoQUJm4K7YZf9kEwQI1/zbRs8gVoc6V
fqCyt2VPc823Cs9gk2XbiCiAQfzDTH93k39OVtaYF8aEEeidEMfpaLTnPOrSLJwZToKMFl25q4Rc
GTLFOTH2GvfUdLo5nq6XSwK6SO2ubrhStjfix0sIB3fKiYtGTGJGlLqkBdpIzd+FG/oEz+XHrDFb
GLhMWGEfthgpAsC/Dign4lNjoFbct4tx9ndPJy2E+Aa7n6JS9re+UqrjpaZcF+yUExoEGdzBeP9l
zuLhru6K0XhLys7wUYkgAsEz7+LTE8plmaqM/tY6hhjBciZRY+PsqXMnKhelyEFyw3TRU0ciQ6IQ
9ARxW1rPnH9fmRgTQtm6V4zti/fsx86yBc+XDzMo+jcqIaY17pSSPuIgQ+2mcihoi4K2FqSZwzhH
rOA194apHVd7HSfMMaydB0G7Al246JpJ1rPiqTHFYclF+ksJZRU8fYPoUXbUe6GOaaooX2ebQLg7
ajspRJwGWdeoqXDHbWr6NuXN7funOY0mSeGqzVJzaxIRUdMYwK4z1tMRTq4I/BEP3s2EcsVppumd
EvP0M513xbmn9baYpWrzZ+lbFIN0K5xqn8BM2bWd37V05pjnXUU99CK5gBd6WsXdg39MvXy0KF6F
XGr0mrbFVaPtynE/pX1dq+k0o+2XKh77b5NnlQV5MjvWAcqLF1dd1Tg/oh91sBuixEQcSChn/RsR
dc5hydQU9gzRKI3cghsnaTQ+Lp76Jvo8uQecgVEVA3KfcKVV6EKJzeTXkFtFlExSxKOyBcYzju5U
6ATyEL853MvnTHilK3qSCZZSDHkytLk6yOihRLFQP+6LhDmdoISo/TNBNufbNM9RovH0uZ8fh+cm
nOAQTJIZFFHI6xuxW60S6oyG+zlGrPM/ygU5QdzEhgEungshNJ2ouMgZ/fCnfaUADhabUZEZEyCw
Q1ghrSfFyVnJyIZN5QZTDBvT0jjUwpqB3yBmeHVRDGwOZpjiIFmFcItxZ0JWlAXQM5rFiIaKdSKn
If4EkZLGZiT1IjMtur1iFkwmuPTnJj10gQop/PbdzUdmi5tVwufRfCaymtZqn6bGcgY+4OeL6bcg
fzqfwz6SvJPIkKC7B+oohbpfqgHB1wWvQEwKkXnRIl2SlgxDp7APNVUCzv5W+g5rC9m/zuOuq60I
Q4p2zMbo6D2QJsaoUSzjiKy4cTZ5WRRtmr3IZu7OX/lswnSVrnKERvifl4w/O/sWvtGOVypctgFF
K6nw8ejAhcBs6K906uHkJE63mm4ojxkLQpwY0wc7Vb2HFUUfoQsdJKhWcF87y+XmK6TrhldkKxJt
BYz3axczbc+R+eUSuoQXuFXXqm8vm+Ljdo1TL3ZjCOK/Btaxq1TLdfxNFS1/cOvwnp4kFY/dZdpx
pZQMKina87g85be+AaskLbk8qRaRitPmlkkhd1JE5X/RaE36Ga0J8K2BYDJmh4+A1GZEi8noVyLN
dqSho14KWmd3+7RsrOOCJ8sdeXh+WJ0xiUuU8+2fvmaG/OKfb3q6inZzlTvPdLOXz/VCpTWjkK43
t/mgB5H1+LrKqvMmf/ZR8WPD8l+SaEYF9sU/j39m3GDYlF4RFVO42ujTqCh6HVuvj0ne72+o/V9t
2X2fPtEWNvyAIa35ZNE3gJ0kbwtQHzrTNEmE2C2yJQ6CTwHJMcgU8VSSdyTIhJaPdfPzL/dF9iOS
GpjBUWCYnadZjGcnFJs+xZNnhAJb72IQllrVeJjjDJtTc20fJ4IKeRN3QGKIX+qFTUXenTIKwtLo
bcaP2uHhHgA+q5w9Bs0fVCV4Tww/vmlZEUKJBKckeVY5JfiBC3TfBN5Ff3PNgqQQRelfle11oiOs
gzYBunl5ub7v4Kek1u87AeAK4bhyQQgmqc5JFHfCHXoXE+bF9q/FD6OKuZIdzCYYipL6AHLU9U41
L5GnhEYDkQK0lLGNnNcVUCBQ58DpiROoU5rYsEXrEEMwwBg10ytuoUawKRTNyrVAZLwVjlUGyEvc
cAC91NfQIKJI0v9HUiBUZVh8x+h+fwOFW/166+MdIkjBRI5SIykB5Pwbx3ZqtDN3WpAlQ8exCUXJ
Xy9JyVjEa2v06WxMu9ysqeS9m/CmyQyVyIfqBB/8UuHZHDe+xNwVf5QG+7PozG/3BgWhyqM3AP3I
JLgLiZZKPOggppARCnJB/KY5JPDkPalKK5QUFEgzCu9jOWsz1e0x7VR9rmWSjeYIZTH+azgPjb0K
u47vT54VOU5ztg2VWjNNOhsdXHNC1e65ZS7mVOb0L9xrbv0dpV5Y3odtF0NlrfO45RGhPzgkw2wF
1/6WLLWhr3pV30f8Da2QsxYKMnFepoiEDk/nYw3cSEXhfEbX2qMZ3A3+eQ6CXoqouoxeJMBI6ev3
ZT0ioqelPZD6BIqBS2ZCuKFSpOwjz5jrOjhCrvpcJGfNtl1Z1mUSyKC7klgIFc1FeFbUgtKaqLor
BM8FmPCE4Oj3UCIzlXzkmVpVp1pUJjRZJ+dumS20EfEl5p+1/2Vi+O/fBVMCllyiySS/FKUAAm2d
qWjtmGNmsDs0Bl7/x4jkF7ks2HIhhGirMY0kXeS/szF+UNcXt7pIWjn3ThNOhxOT+p+MfTA+mDNR
lzBA/naqIRfDjIcW5glqegsvEtIOWS9THY1NlUNOBWZ/ZOKhwcZDF5TjLQgZtCh9Sz5+xkk6ucxS
dYDqpf3XPXikmB0ZQd3TxjlyhVEYSHPNa3vcijAgtQFbTBvNCJv5fQdY7RAxaZLy3wxNEWPw/PJv
7xS2GZZ8Kf1jIP8XT4QuHxasjT1R30qNUWf1JjaDVn6bbjs/6B4bpZm9THec+SMZQ/mokU8F+a7C
a4OEce1aCitQjEem4WcbY710gDfF5I7gmSpyZmosQR8VpanI6S4ET165Z0ANIz5zGY2TqK3ZoE7+
JGzB2M8DpYam2KTenyEZgw/gmudTq+i2EkCPWCRk6M8xzmlhU4r+/X699xkQb9tCaCGTg1NJZeco
+ZtxO0jIUwJuJu7onYgUKDhsQS5CdgS1ViOW0VP575Yuo9P/1HNyp96/JTaNR5i66isFNrHhkwc7
fHmDc40mPgaPvFnaErX8WC2MoCLRu+mUx8eAI8E6x3ZYDhd3Jq9fXINHm3p2CwrHrP5EdKtFRlPX
/ZherakJUYC74m8/KljZJMaQeg5Jw1hatlDFVlF2StncJszI6uLUH/NM/w5MdShiAn1ph5NHP0P6
Al97Q8thfP6IjHNRygdnBN+vWHjM1eonWPM2gE32PMUWLgQYgN/uIOM6kwQSRlT6KOfTy9lNP+HS
WstHqHFD9lEYiIY5NpFxHdJg/RIgomt3AziruG1Ntnsc/BOsRrjd0HWzGWRosas2unQnrE3D7KEh
fyp2Av6kibCkvaW3H18bx9rs25Q0JPNCj63bCL1+g/m2o4FesCV+x2mPpEujrWBvYzUJ3gjBLsdT
kkYT9pL+Kqd+Cf1yA1Bd1NWUg9Kn2hp6yCHXK9HSYttAmzSjDHJuJ5oE6FRtE4LgQY81gXpyps4G
PELWub5zwsmzmZ6tXvM7oUZQXy0l7nhmknk1j75ZFFalGmdGSaS6ukrYsmx90Q7eh4xPaw3/RiFF
S9syXVL4bQ4VxTrLKHIkpejkmByMcKQzAQSm6czFsgbPAtsrfcEl1fU3rkrekbQfsKXZBwrQMLT3
0Grq7Movz3ULFVvnxZYdGhv51BRMyFvfAkHBZiNjNld3HGnYPLO9F+RIJMfjcmpZaz3bkQ4Rrm8z
tRCEWgqtOZpAdm/Wjt3vieCQfU7gPc3gboRogw4iPUFay8DhZb4FHqZUthzMMexouV7/PHDDmVIs
Nd8Hg62zy0DTFLRzBR4bJDo7auyjt0BEqZGqFJTPE2Cs900f8FzphVgVka22NQITDTzSayf8oSTb
p104dvLFP3+ohUst8jFFaTTKpE/5erzs+8kssQqD1ZnQOuxIi7zsbx1YrEVnR0VsS4+Z7zU/LTiZ
knK3uvIkXW0MORQ0WVJuU3qWMsILlkUb2VY0twyQ3DrxamNLAZewhoh9iVLrJKyt9pyoFxvD2ZTl
3w9W88zzcRcR9tGSKfOoU3IG7Iz7bFdi+w1VgTRPFHMFX6d1BEts2H7n/DfhUhvMHNsXK6yn2LWB
gGkFHkhZM+1pFBHPwWGtMtZoiC/EYh4g5z/ecAqkVZuUOoa6hIyzMJ1JzVdWAd1DortODnGUCoIU
jEBPzvOt8hgpGGSTOTwvCUn2DSXa5AoE//vMIjHe5aNwKPw1VmJUnd7kBjrs+VN2SyKRwX+PqYpF
GbIvCJCeETOlVC4uMJUto35Ws+Tt8jDUU2x0ritHOPU46Z/NpIP9NMiECvLnaAeU2dB4ccl66+0l
JiXti6VyvzQ3Xn7G/2ek0/Qoz5e8vau0gL3vUmXaekAB4Acb1PiQX6c6bZ/bqCYj7Tdm5SX9PFf9
EnDizd80oVIUo7cWrQFoGzA/AbFPwdhZyHdUp5J7CvnZLNSsJGib5sGzmOTkVC2dnC9sH0sYQJZu
YvfJETcWtXPx77qLJsjmR9f/S1DEs3zaAJica8fNZYDy7OMiL25At3ju7RMF9xFc8wrfX/J84X2m
7eenZ3zuqcTa3NyRLqMSMPr63XW7fT21NEqh80JDclsA8KDz6P1e+E7Lpufj8Z+x0teCiTp3WqYy
lZ+KrqYq8ecP7/JPq1rd8PKgaJ+RTl/jBenCIg7ceOqqGRHwKenm3SFGe+YLGsUvQ3EgCpi1+pDP
uaBctj8dpDZtzYlTPYgO09uy2LDfbrY6HKHtM/rwKxefh/h4/n74pFAFe13Bw7Z2NbMZvAIDf+29
WhVxjUMc3DKmzJeZFqQTxzR3yuZbxj5qV4c//VUBNOUH+IQIc/p1Xix+4EkTdH9nSLOiQKjR+iE4
li0evcnfWWb7xgpkxGI5B8ijh4sgoEGAiX0OphZwRTkYp+S2WbfIKvCAu99AyT58wSH95VOfarLw
ft4l9XzDXTWwrhyb0iG/TYjVkwmD8Mc17x5ALeoo7rdz7sX+Jd4Jk1fz4DNVP3ywLvRZglykDteT
+7RoYfxS9UTviB3V/1O1i8XGckVKkkozp9krB4w6BF7n6W+oFVIuMos/ht1ymnv3pSiD9KgGnITp
bjxqGQ6eQzClWW9ZGOO9QTSNV7qEUJNpnBmV0FZhaRbPv3COPr8K3Vq2RvodCmoi/lJ+0aqSQCoU
ZP3A4o2+AHISDpJBP5oh1xJuF7054UkqAb+euAJ0t+v+PcCh+XESxLN056jLnX2DGNsycpwAIK2e
GKoK6MJ12P7mFOJE3BU/6d15i2M06jLuXp3Q51lFoDdZJHj7SEa2+7BmEFtMSuvL1D+Qgl9bbsYg
i6D70+PVS5Kig1UXomUZXHp/FA0ontZL9o3GAWXwoAvhBgzC31u7cfgJkcgpFy54RRORkc4MG1OI
Bt/1JCB9lJbt7+X5cS+fRhQnTW+sgIglPi3BzSAknRkKTjM6f7ZgRzv0gzd7IdIIhelD6fA+t0iK
2nbN+CLCvOmpLDPrqDvZBKFKL/5deFd61WVgnm7JLNNUjAzPzAXsqEWwR9VhsMRdhgNdyAE8UXAa
W2OA2ij9zFhoBMtXY9SQEu1ohy04Erhn2jEu4K01R8m/Gf0PEguOMHLceKVeoTcv9o40vp0Q9hGs
GlnvwFaf0gGYE6rPtM/2kSWy1ch9icnHVeJYJ+LMNFbs83qRiC1Sq9/6pTT9s3ZHfmORV8eDfvXa
Gak8Su3cj+FKuEVVOm4VuWIhxekJZ/L2vPBtDzYzhzDX7C8dSh5G1/OBydLUzCTlbeOZmjPa3xKP
vOiD5JznYSNBJZa/AC8Wub4O9vwjmKSG3j2Y2yG/2qE+VjMkZdWKSyRWqFA7DiX7g9igQ2TZ/TRR
FEhPiWyey0MiXT0xjAziXsKDKa2XzHhy37lsvv+jsSTmZYshxz8zRnvj2PQeEBGRbo+Hb0hr7jR1
UUHL7IjqpsXA6RWNROpQtRnecjTTEOFvPhwVOH98se7gcokyutsspiR7UZLphyV6AkjD6KU9u7Ag
JCLJLIFf6zVx9af1THuc+yFeqAI/Q2I3RlqXc3Ow3HSRQKWpzoSv98wJwWCCNFcI6nkGgkfcE6IE
wAoTNaWHJhvWSArbx4iPpiApY2uRRCkeJsv+HEBkqYpNVOlL9EtsDPI7/iWMI7DzQgloB8haxYXo
rk0wr5I1BfgEwh0OAWo/wBmm8kSToIQ0JvTbwa8NQJvV//B/+llbh9zhdsLTrSZiOTVz0QZoMaZu
8s/GMfvKYIcC7RfRA158OkxNvbG/MGZwAtoaMurvLSDmsFIQTHDzWxvabYtr+w8QEnGnNOx9doUa
ngLH19Y2++uDo2MfbiEeP67hFpj9qdAkxS8Pur+mz8ZuKGYmckKe6gFk8rz8cwRVrqeFXiR4Wqqu
pzjn4T8YmTdsyAk7BOht4u9T9P1kE2YcvwEeo+vWnJW1XXHQ7KFhtqBVH1dDytSIuK5vlOGpF28A
id8RtjRurgTSQ/b2IEXv7o6fWgwiBC0wrSgOlg1avE4Z2hQlhXjGIh2+RKmgxv7tD6lH4uMOBqc2
5MnaSHSU1+BO6FAPsUn9r8unoLon/c9N6MOnWtAUKf+YMtWyuHNVtqOIh+JFBkzMg42/MmnF49ML
r6mrWn5kbbo73YZI2b5ciAf9VSsoktl5YXZ6DmFGO/z141pXH/RP+7Q3sleZhQMGfFIwBqRvhUS8
+GV/3z9m6zmZQWOqxKMVjAgL8+eNkKP4d2kjODA754Ddtfsom1++1PxyEFTwT6GXg2MYXCdT+8pj
kvzoCDKv5Z+uaiX3ka9RCooBCOR7OAoAyQewGsV7CJkYENcqyASvX060Ohh3aXEc+RsVz6o8e5wR
33Rc2cAn98xXZHQMBk9ZpzYOPQ+rf4pM5LZzyJT8k0igBw4RIiUu+tH0Yjb3kte4efx1aX4xehBx
O5PUCnId58HCCazvOY2fJPIVTRKnG3a3bLTvlSJfhwaxN6kV6IYSvh88RIptV7zgwtaPe1o71UR2
WwjzCJKy6b6p25281Y9tK8Fku/BjnrF9xKwQ9mPMm8bvWiSXGsmEEt20ipQ6pb9MnbrqdCzvgjgE
E4D8s+6tCweBpz29Llr+BVqXXPK2MpYdDuXS/TLyMgrkZP3LTvl+AG2kQ3n4b0H8QrXfa94pWBDc
Dm3t8vEtK33/dQbdpbiu2LZVhXV/L6dCUZFx2LTTsMM1XfTJH1ij/cLCW2KBjDCpCPTSBVNupEu4
xjetEQ8Rznv4PZ7q2zqrEYTQDt6+2Wsg1Uwz4hEXPKbUWBTgtq9iFKzNY5wTNINQoF77CWLiBUca
VrsIJvDIdjZIMDU9PZtxkX2W3/4vPwyWCLKiBI0n16wvNhzgCWYi7nJtBtb9LRCnOXRzkz8FlzJG
vr5GtiFvaVK6f9zwBSxRx4iVs3s/lR154AXz5K66Fp0aLwM4EVxGwz16CAPBzOjM28wW4rA4QnfC
x99cC4JwCyTVZHB5vYNB2FDAQys8hWOiq12IUQHRk/gdJJyJh97tVR6cmsqsqO6AcjeZEc7Ler7T
Mfg9xPMNMaqGJ8dXVrfbOSd/pCGY6T+8T3F2GnC+2EAl+UjAgwsQ1FwKvkCMOGgcC+d1+9hsCdw4
v5SixqhOC9aMqrDkC6IzZI1sWFCdc6NNHTEHE/Gs0TTrzvTuwnSuMPyJTwOwXEdcXFpOHBr6Al07
J4vhvJ+HIajIIHK2bgutRl5nL3v33h33JsE9uptn6x6316WlLwiNEGmCGd0mxd3bYo/XBMuLih1d
1Jiovk4ovhKs79XgoTKlNYaJ9qjctwRF8LioQwCBToJf5rSG7Bg1HgpVVGyDlokxny9/kn90X2gf
kwFYQokXuqLrXDdm8E7CHgYhwP2unJoZGh4vo0uaIq0b2bJBY95/6peFLulxVcrH7UZqfnQzsW+l
46OFcW5fWFtB0/kc6CjeWq7rMMnrXVsntGMj9XPxpbrsUW10dzne2gicwTeBiAokqNs5J8N3volX
3rfQVREu1HGnvaKQS8htHCjDY9xpuToQwg5dAMKZRwdJAJ/fw07mcmNdoZ46ihE5KNwk4fbfrY6u
krkRmWWOTzgyegmKO49Osrva26o61MG2esnuWCqym7Gj7LLNfT5dkE+R6CfORKgV7uSnyRDgJU5u
1uIIKVhyRzO1j3CN4NpjyORyI8zHgEiWY0S0O7QKDgSzvSwmGeNzt3gy5+44uW9Y5tn3Q5BofN7m
HNn0E4TcxngjUhtduOreUihY8/EvCi9nj4+yzkCt6fzadw8LXD0//z5m2gWdwzBw6ywQqKS6h8fj
/0kAl4uwmIklAUfnZvVZvWlBAC6oeqr0dStS8NRhBAh1BlfLygvUAmlmMq6RNJLwZLKGhc0egG8k
XlqOHbxm6YHNKfWcvWXeAXXjkiJeMqsMA7sZ0g8GsA2d+YYlIO/C/wIfpAiB4KsWE/hDfa5gJolL
9a4lnAfqDKrVFNp5z3IEn/yEdJ4jX3S6QMEdYCiZVbIzmnZNsH+iRHTbzJHmlOre2lQ0lRG2+WTs
yxKSZVYPG+qQe9pW3mMclRsgQWBneo8+qOZbbQ6b6PQuU8+IPp5vwH7jxHnCDjeBLWCFLJLcZR6e
pBHLL/opC92uc9HuIjiZFNAdnJBS9P0xrTDiRZFVx5PR06VRfw8SrhJElPQMkQjHcYfNMKtO61cK
i4Wt6RsRDv/KuWO9Mqv5EwnQYzmrOVP80dIpqDrDAQv5BKzcyHizj/hbbqONNkKjSOp6OFKjBWxG
8JytjS7whGhAWYQsA3lGjo9gwtImLkx0+5wLMRq6+KOTx498Z169CuiV6LG7MsWF+81NHl9MuPZx
IrqCB12Y7AdGRCckRf7SEOzesjSdrEU2CAfWAMeW8/5WTvQb3UEtEB75qbGZKZZzmy0ovUie0PsB
3xdF5oqRdnJ937fPYbD9nBaX7bQ0iEhqa4a1B/WBPEz3ILPF1pEVoOlY+l4+CjZwVhwOimb0gt7w
uUVqVIphnE753dZkde8SXExSpW1myanmKAnS48WXeK8jy4KsUFIs8bxWcQ5w+FLVv6YZnESYnU0C
MvZnlzuXxXDFyCcrLgiYCdFy9ZwypPlgrxMFWWE5t8TOOxELdNk6Fi2/Co+fca8MU9wkiyrCDWZf
mcO4SQtnvDZ38w5o/U/MyNUUxhdvzevOzry7QHuBAG9xfiblT0WlZK3gfbEoJhPM4Ms+g4NP8Cgi
5uQf85nNCHkKO8shmT2hoKVSeu4f3khv/LZ30NnXkB8uFE6gXHXA0y0nWT1z1VFJWX7YwgVv61RV
EYiYLFGc0DHz97s2xcCYJhmn7oNvesJjMZAe6sH4867pdSzMDhVx3x2IY3fzNw8TZtOwPPWA2exU
QeN9SZvUkKL8u2zatiryUBd77oI94V05rfNHRRCjb37RX+xk44jRVKuPd5jTVDYtHxy7BFqBZykb
J/PFjw4L6alSPiFVU5vB1tnM8ueolj+iZWYO8eScvGjTqKwhkIx4b1lb6TeeMTFBkBWh5Oe9YW4A
vH3a4OvIJuc6PZPgrkf1J1R/M+R/FBAzvmy84CCXvpD3MlXy2isnfkGE+exrI5yHWDr5qxbJX+gp
cPjzMWIu/canIHohzKBrlwFw9IvdKTlHtGwe5MOQo15wqALJq7KHyCLPyVl5N10HeSrtwBZXBZpn
Dcwovv/qyjb5ui+AhSMYH3BtO5WrMH/1FHznk4/ShcS2yxlv85HnFZ1YfbkZysVXYvszp7EjsF4B
LDtdiO4kgWwfFC7dXrWTUit1raxVjyQifsXIdogYUa73dpyvrVMz+UC9ky2KguE4dFve/wGWSIT6
F52AEI9mnRFUvNQ3zzmI/Qucj89LAkhISz2pZEOqR9flf8ouY/HKgQGHhvCzElO1m1Ojx7LfwuQk
pn8nLJ6kckVyMz3GJACHgFHCRXTJVpnTeeF0sQr12zc8EdZ+uY7zC69acmZ2PccFnvHQ6BCfNLHz
2MJXDDp5Cb2Qc9D09vFFBxRIc+L+9R2GvkA0JzkxKD79WJTOiDbFhGxWx4lcRqYYk9E4T+U+37k9
Ogo2BiEb0/vrQB3bNirnptGskPy0yDyOn8L6e+gGch7l1SPMTGhQl3N03jIrKNkOFGzdttasXdQK
RTGbrsWRbiQEbZecN2u2JjQ2hLtdKR+qU1Jxm9TLK3ThvMdYFBqbGivx1W+e3FR33INV59RXPxFS
8Q9V8I3uNHxvNYlYTZ4FMZ6SvTFZHOxuw+xwFd8GLTF/uwGvt367X1fH1cl8WsRn33O9K4rff2sW
DnZrnsQBZJoFME0DikV6Px0yoG+6PvtgWkMvnKbywjIEI8FmY2v4l7cZ1SjSBYhfS+mRflCYFr13
tRRfVXQFPDYLyZFS0MFBBklbxzn0m2tVYE6n7traeaEV5L+m07E7c8bknYdMCG7HpWLopjkXsbF1
UoinGJMB2yo16FCQqtkBwjzWAc+NpYH4ppp0HBagbWZ4gT1ylOoRcuuAqp8lgULSFi37UmsRpzTj
f21v5YNHMUrcYQfimsBdai481kEbFd7/aeNEmyDGef8LgRAIcqSJdMtE9UMLniRG2L7aakSMJd2r
VBvulmXxGz96FuuR7KEq3bRoZvHmle31noF9na9hzladuQY/lxig0kWBacRhiVR9xLNVHXiM52nu
rNkJx8yfQmGxo8kVZk+TglWjAZa75Cpc4bRXzZPU4wQEjQdI2hj2o4csfk3xUUg8rBy9ImGhoc0v
5U8AbaDLGTnkw8jG+A96yyqqAImac1jxRxGO75aLVz5ST5bqbkLwUy+kenSFmd2c02Xbvgxd2cvL
w+GLcPy/tAG3wGNWpc3SKV7NYMCnVzTTF+g6++HZwX92FmCkxvdZKtFKsRTwGtPVIIOHqfcra5wo
VZgU+qQU/vK1lodM0k5rOIsyjIhug2Zx6Ja+xdDN9Sv4mRnWOEBoox9guBew/q+vu15gZlzH+68/
62qsjDuK5Uyo2NCMS2ODAXC0MlyLEKS5sncuJedGqS05Lg5vBlftZooxd98Lh74nahlURkWPpzRY
G+4odNcv2QSIukWb0JPGFC5WAaLDbfdY0l1OF12N6NZcQ1x2u3MVLb0VQdfZUxWOuJAud19CbHQm
3+zcf6jHaBE0O6dIPXNlVg9geP3pzGexFBXG+sm9fCaR3NF0HgeVYRpEu3GRglILSLASglCXhU2A
Thy32AP9jNIxHXD7QWj12+ckfWdBTGapQOH83c0SldTtXpROiVf7pKEq5xKsIH9OC97RS2HEpOdA
pgxCsvqzG4hy+ssZobicVwqhQHVG+bdZ+0vplZraqFggRnG0InPaxkJCEH6OVnfojTEbJGk4LnFH
8+23FuyebFuDnWdfZLW5Dhnhax2r1DalMmv2m4VdingCRXhI3gz8bts9ufVuyjyu7XQnY0sJAEoU
7p6iu57H4CLVLWT9tiQTftpKUjiTWfA+DdBnKI/v1jvyCWit/HflpI1IjC+WwJTpDoYCYwLGavXt
hpzKJ3v9LG06K0+HEw/FNO0BK39m6rLBSxuGuQIn1+iW1bi9N5m54VXOJii8y8+vikM2ordeiIfn
AFjgZKykVoF/DIEXjdjgk3xk6NmbFTEleWFaM6ZcKhhpIqgRJNfLue5eJh/NbmyO7+maJeobd2ka
EWa38yhp3wU2b5MjVKuEI/RtTFJiOTTUy8pJ9ZxgTdU9xlhfNGotajz64FyofHHBcKaCj3b3pRrw
eLkTN5Mhx2TI6140WxbiESFJhDIwKCSbTwQCZ1iGiUNyuN2PhlOiNgV5rf4V1fTqEP7ooxByIoHV
tCk+I6D42fKDTG17EX0NtVihQ76ti3uVSsmsnlGKhoThuQRkRgJTBfynlg7WVwoIvaymrNQCJ593
aZ8n9Ivpwp2LK8lT8PZsYkB73oDcakQ9jjigOszDK9+/IRFiivq0wxW2ph3pRr7sBhpCtw8Wbmw2
z8UtHwbIDF1dRyKbdtoImLt2WVpWnJHkmCVv2YLYgIbCMwGIwmsrs/gEF+SvGmKF2PXIUo0ZujgB
V4sgDECKPr8UD4ydka4R2XqsorfqlkT1I3Y399KuGoL0AeFLRiI+1emxkeV3hBCPO98Ql0pohlKS
7V+A3i9F0somNkE0OuxrmOvR9oXAQfzBLNJs/CkwI+Bx74FKX06cr5CFiB0Zt8KaXJxccJ+D2pOl
Ta5GeRd4mCca4Kx8a2P22Q04Cuucc+ond716oN+LN7/zqnGUjalCIZkq7Ku8HN9W+dnoeihgvpTk
bhVdiAlfinG4IBvZhxvIuoc6pJoumPNfZYn1WkpmqOUS3PYpDl9/JlFf8Y5WYA9dT2X7HsL/weoV
vBcDLC8H6dYg3bodrsUd+ll1q1x1tQe9/hDiBa39jZfE+IRfAY4vZLLyikZkS9hFqWk5TaR3ryrY
aL/DolSnumW1G3MozJrHbPdnM1D8AhX8rXjIT2/+DUrqE5qqz/Nww0riRwRubY3eD9Q9Nt1MPW1i
b71Dcs5I1vREY+BKXNyIuOQ7ByDBWb7VDVn5eJEQXd0fWlIwe4Mp5uB2EbCazsWLMT9xH5nSpuGy
vQq7q+gljhBgNxPuRFz5pH7/YHVpm/xc4VYGqQyCqoEdT6fVPKz38iXjrM7KNW0jLPdf7mDdYulL
iHAr8Qz7g/e6nq2GbGi0VI3lKs3xh7NIrRYBQm3t/xOuEF2+7LWWLedUEyOZhArYX9LlyWYPIg9u
UEKPIKKwO7SjC7nWKHUQKmwLe6fIISBjqeoWZ7u8pocW6OW5frb8hWq0+yGXDaxRKYbMb74suuQw
jtJnozbIgitAr3MYu5BWcurJ+LYELbXbK6YAf+5U8FuUL3ENdYPNcVhljFFKhmdsZ5a7ed+g9wyt
Yd3E57pCaNrd8kOKZJzMsFycquhJLUpFBX9e7W6iknZEoYeugw0Ad7BGq+PvpsuJ4nK7WMSqa4/M
UaCX6KoQ9tmuvCgNMA8ssjHeoVS9x3oSnBH/qgj9Z4LWqfDPlDFTJUmjzTE85oUkLUBTlTG4/xP0
0ERb2MP5zDcBFa1UIPw9WZtaucBytQZuL+PmBYvbRZo0C61xHV47tiQc9BlZfILGSdxAtlmSKQrk
T9NlCmMVNvXXx/n3fZ4sQg3tBbmW3r2t05YDTdK4pN90oONNTK+nBxSp4fiF3yrgQXRSXsBfETiv
eGNsTdQ5tJ3BSTnAEPLdEAlEOW3Y0GdhJMegAe5zYtSVYX+RO6AUa87WwLd6Wo0eegh91OeMBGA5
EqsvZg7j4zuiB5HWj2ZxN5mFuH90Bs1GxlBR9at+HExj8nc+52NRPol2oaarR/yTWyCXQigs+w1u
4Ao0isQVm5PK31TQXe5eVWag1oPIx/zj5pJm5IOk4RfVl50C1IMOFz7nC7GcYecVCpj253o4o3da
T7oz+lxQ0/+Avxc6EjcSTEY0n9lZL76CFpYAh30z2s/1hQdeiEOQiyEKiAwEPxH1SZGfypnV86ZV
VMNh7Zzlhk/SiY7Zv0NPvlISCKxUTsEYE5wys4N1jwJSLxvhZHsun1MXLMpk+4pLZPkcNGIThWFs
rW7D6+EuuJB9NaNasmwTcCPWCWTOH99Php+5ZGLRRr4Bm/XYHEBr5aCTkhEx+kGJTvGUkRfp+W3p
WHOcdyy14YIGT3v+BMgkco08/n+V7HSOY/s3w5Dg7uX/qmxjXsgF8Nq2Cd5eh9udNp66P/xrSOvQ
mPq8Gvh4/KTwM1AaoP0+IhfUU5Ap64SE08GiX3HSL22DjypMVlLzE5BAsb+DpWOZM2dBZiqrpDBr
Z0OoDypc66JnArwRh+7AtV3TYkXrdsePGALPs7EPaasaRSho3ZEWPwXwfws9rFGVx+1mHc4Cu8Ly
rYLQKqWNv310IXK6oPyDlkpRCa712sJV6Y7fvKLc1oq2pken43GOA5BP+QIar4GABN4b2dHtFcKm
ISo0KBEo7zxGWTP4A+srieMW2rOicFP/5xoYbixDFfs5tma4kaVFzfUj26VFy7FChL4x+XoKrMYm
/RRjKhJpkBMkASEdC6pTu8y5Puu5sn/sURA9fn4gz4hQggvDkSmteW8sbLErcul7WHy5+4m7MEcV
xPoUHv+tnIWqGCAvqp8Z1rErID/upXO7JWUxxMITV7YoZcqC15Q1pjMv1wqWoq87nZsuRILpBuj8
/Dq9XhmHd9FtkYAFw4w38taTmMs5Q1lpA3f/vgyAzGReXJvewzAuD87mAZfmuee5FYIXU0lKbwV/
57rySU0HVRUCqlMdXikWOD+yWanwuLQwev73nwGDrqEN67lS4+KY5RLverOPK0cFDC5a/0kPJO2Z
bDrneNXIAWvaZrlmDG9+OxHBFlqsUO8GLm2l0s8mooZKj6ArrhtVqjfjGBc/To1lBwqnv6jgwoFS
36gHchom+MR9ybxLYg82Kvq3qGwWEYZoyGMeE3di066rCfyK28INLSKhIheJsu2cTBm3RU40xldF
1TFF/awPKYb44y20R6NaH3DVSK36ZVYXJluwEQTSxvF5voNPj1vIIJ9WalmfGzQE4600SFqBPwvD
FdUvWv6rY8YGUreqGfE7w5ory21UbBA1GGHaa2wz16YG7xYYd1rcfNIaCZ2+b45cXI7iOMH6FoNl
D0GMGm/ZPUiD1/Zfl1g2QlMY62YSmh3gVN0nmvFkFBsP+PvIDDRlfvDQM4wviYytbBRfXBXQJXmj
hWRGnFDcTIWqeGLDGDggdv/o55D89s9YO09x7vGPI0WlPg0ac+psfd7+biLif0nU+qUos8GRwrWM
M+nMyKd8D86NkcD3VWxGiodtBMP3SS7D/UbdeYOG2ae1C6IguWZmex5snj2CGXN+zqHfA9pbY2J2
eoTcCwaxU4gpxqrRGbsAGYbO0aN7V9B5avM9TbVZlRqfJeKHpz20ZCME5qZpcAnRaQq2lS0jkPdF
M5JPcrLkWwz32hckQCsWulyZld3w1G9CDBoY4zjr4wfN7bRhUFYaMONYyERVt4ZH7c2dkjzs6R/j
SWil/ImDZmKytVtPPuulwIjA+3FzXRFx8JCUyywdGwKvZmVB65Ty2+QyBSfQRw6aF5yZUKBMYJJS
hlKbUdEic/NMQIwa3D8WpoJcB5Xqo/Ky45lpBaZ099FOSiUBnenmsqkhNVFsyoeDOx/9KwZgNygF
2LpsLcyKiXguACbT0JMb1YoF7wvtVBePkilxwF+Lxfas08MTawy70/h2+SGj/KEn/6rtNL1BxTbu
a+plITws3OqYN5fPo2XRzlA2oTyk1fmBtm2k9oDxw33GKrOQVmbMBRIiczkuudKcAZodzJR16I1Z
qgLOeM3vAF5QilRGJ/p4pu/fWk+hpEIugyIjki4fJ/x0U6XZGcp/R7KtPOLj4qE3SLnWzyrk2/FC
lvDpn6oYgM7h17dZa4Cyq47o78DphYaBFN4jaCPOK5Ei+yM2eXYftH0S3SACGcTXRyR/QRgie0uy
HS+5ZEoL5PdE2dkoo+1Jv7JFajZgvwsEict2PJ9inA7ifFNNh6EBB06IPN4B3MqsyhQTUEk2TIf+
uH3vDQm843vFxe0+3P95U1hWAer6bzdl+mFF8iPM/Q+Hf+FJicW2eXGXka5U0jf91UT8nZ7wZiJ3
MhKARWd8LAAJG8L4pVNCB3wF54oDYj3JKWYgfyiYVajGlGvS1wtc5i2mJS8nBaCm5OAPet7J0X2E
Hysnn8yYun8ZpM6WMB/5zqQWpsyh6mQuNp8EAhIECgwtGBfm2198Fv8PUVHqU19KZoEsqQm1t6NX
JCL3ZHz7w2RR6OeglBuUifFOfW06Ge0thpv9kmT+tQbie1j03YOC/xb0MItTSZV5vy7i0xhh1pM8
eaH5LLDo6xbW+b45qRr2EepKVXvHqZA9bOC4dOMoxQ2v6jrOfW5WgoWYytyE/tZl/0ztJulh4TRx
tbllcd5FP+q0TSznKujWLH1PEe5vuICwAZfQIiayoBxlhsfBXb62P3xPLyIlStC0liu2/KRHUwaT
Z3H9WaQcnLLlCIkxHdPppGGVnyVm8Wu3TdM/DbwwOnZssfrhwjr5nU8AOSPfsNuHZwFfBKjk/O/T
zk/qQ1n0ppwUCPX5BN0RJkxK9VqUJmgkKxbhKGEZQajLQzsJmIALG74aNER4uPhJOx6ZRBLEU+Sj
6fQsSMHunj3rgsTljPZojO18Vgg/mYIyOaAnnhkfuIcsLglwRbS5czLu0VhY/XEuSSqWW3LlNEYU
BNsKNVbO+/vYORvdsBHaiGH3AgH8g1k3aUD3QRuipzM3hrpTN8js4RsdoOUKybOxFE2EqQvhQcWc
STAskHZcYdCqfA3uG6+7S4GPifnVDphecKtnDYZ2dUhLuT5y+3+lEZ03f4wWtkYtELytawjyGA/v
GPJXJOz89oCjQsZ9Xl2tmlL+QOJMzzsjGDpIEfpkx8S3SAEn+kWCPyg5h9hh1ahApDJHSzXQiwPu
YlFohR7dK8P8DiLSOQygrmSP+nZ/C+WRtEazEW4rZxzLidYDnK9iXtjoLJN8zyU6gHkV1LKnvhtt
UQaI4/YeSqoyW91b60UHOYINr4EkhYz7MYuNY7jp3D5GUXJfT6oddfgay6/2yHLhmHZeiC3jqxmT
7KiE+PmHdYd2ZYThgpVngMfy/VrJSyJ8uOBuUeS0wZEo5QwGB9iHWVWvCPjUUm8eAgoTWEO7Go7U
EUQ2cpxpfP6yZM3myud5EW/e3rssBjRNCo7f9qYaw+CBPRqYldQzXRfnpbCHcrBQlkB3YL0wJLVy
4yYhfc1keIj/6wDwYoZi59JrGC9gYO12st/h4v4yq4uy57DhowgbsSzeZJnE87ihqygpqYi7g70w
paMRF+YOQB6NxwBZt4qP40uAo8kYYZ3xY4cn8DZVykw6XFfw2lxYyF6uDy/GcWzOgZlmoFqlxfhh
wY8WNfvDXrd33gS12Oc1DJtntEg5WqUIsRl/opoPp+gupiwTAeSOl+DFgPAAQZS4JcDk7iVw52wI
PHfOOlhqHPGh1LTMiRLGe3OBU5EOrias2EVg88Iq6VNAuccqGJ4gii43vSggCNUocks2kOh2DKbJ
DYCgRSgzyY1vov2y/Ms+NX2McHg6vxLTVnFLK7x0xlb2qKhXYM9//zyJPJdFugek6rkdEH8ETSVK
8SF6rfShDJXC4LDjXW//EqrsdF4eOrbUV8gzcoyT3ioUstO+6cNeQKbyUkznOeA5jpd0AzlblsAd
9rec4vZMx565IdDNdK8xO/NTkKx/RWu8MEjsCaD4T1szaP/O8FXBLbNbjeI/gqzqzQ1WNdi4rFCh
GGPDCkiICUXcNm2ov6K5+TzOSP/RLM3Hpk7kr7cKO/YtMTM5ZXvmIv7mados8R0hdGYjWiOygGVw
nWFRAhoHQuJk0vU+7X/rO4UsrRk3rPryn08JwSQsy6T2DeVvEAndGziteOoJJAYWVYPWgkGYR5Vs
2cFn5NTxULODfa91yaMTDNOxEPDC8Wpl/lolrYDi+bEGSXVWgKAeIU8vnBCamtvLNl050v8pbTCt
EjuX1+eMWzApRPcy0ZZj2mqvqqt7HGwtYVkCGRbOwZTLH60a21WIkN+UEloD+3CES7Ttdg6XzL+X
E2hie1+R20cacA8P3aDyqLMkfyDuuCcLkwcrTQf737LSNEXjs+nPEnwDGpBErmkK5QsmmRVaj4Yj
eIZ6dWCjdk+BDJzf24PCdzXZLCzFiElbfIkC2TSfdmZyMnBjB+CwJDtRrwS6m1UKxwkPdy6a/VTL
dasyPrhjgn1odYbDot5IENh3+qxefUOBv0u+19WRxtQfLDNdXTILWd4HrFZTnFGqV5KASuqsPquf
RXJtBsQh7E5bgd7bIJyKtiyvAOW5CN5oP2Nk8alv2A9KDjCtHupWcmn92QZ165HbJlyhXxebn9BQ
5TlNOYXAqAQ4CnQE4NSyZAYB6NAuJ6bzKKFtONE46/EPVQ8tjhqhkkOtwpNCCGoXldrKGdDowpjh
lsUEqjbN1+QudmcqAoFiN+Klt3JDZsOj8ZxGePjR0+4RZZe5hojQTBd6ZME1px7VoC0ZxFwO9BF9
O3Me3xa+sVvb4ZZtArehQvE3UR5HS5olusZlPBmW1q4QaFRWDJuK4LTaeKCkgwoPj4k8EnDXx64S
H30V2L1047+88qUwR7y8v2vAiwrI9+JIVG9hmjkm/9k0QChqFowM2MGXUhg1gAnb7JrIHw8sP/GY
mxqmQMCvKvullwPDHfbzX1RVEuRamB4UBGQvvYZiYHrVOoJypDqjr4PLBE/QUi5mOGAROHEwU9CQ
s0a21jpICZxoiCHgpynswmTmPj5g5LPG8+Vb+W1l3B+oBrO13sNlBYhSNGrB4a/lQg5fUQF6aWso
QWJo3+s81e9LzGr1IBaCsOrcM+b90bKuC+GulKXUszkX8GZ7vOYDdj5otas1f93MV60EkCv+UbVH
DgffIwOdm6dZIQrK90q+jXhtgZ3ObYkRZJJfoEUI3appVkcLDf4NaUPuxS/b3b8diWnm+XhExMp+
IdyDxfdO5L2WAD+3kTjTfaNmMPT5lR+oa1VYbJaNI2Fp48xbS2o9uVIuSSK2Qwdm8hvnM3bMJi7D
+Qaw5gFpgrG6oqmySrj/zTbFdh59hlvQ8QB3CHhIxETUEJHcnLt8j03J6GKp/qoi8z/wVgAFXwKh
RzfIuQVZXbWW1BWHAPN+9wswmEgjvuJaUSNFLaGQ7Qb+5WL6oLuhiUTFra6p9t3mKnC3Lu/GLvkY
2jj7QUPuVG9q08f2WGswyCRjr3tHmlZetzI6h03apRZBTyvjxe1h+Dlf66VYb9FzbEmCYmxUvSZn
/eAe0HY/lIEUdQwEKshq5OJN5kWrKkRK7QgM5ceA7piJ44lXlxMSwmn9Rlh3PAjk9DVoITkFwRk7
Grlnw5jpBB+jQmPgSykwlGy2bAMU3X3aNa3jach6hoMY7XkD2iY1xUxl5yGL06kycstaJaFMQc6S
679edT36QDmzd+3narVBQifXLRW/uwj9+p5yIpEBgqcgouBVE2ad5Q+63RM7yqVraqwf0H+Snkqg
ITVNoN6KHxeYivY8UP8neBbBMXyz+N+2cT+3zxCIrSK/GKKlI0jAA36K799TUyXDc8x7YhDUYfc1
xOvOgY1GDZUVAeZ2ZCh2fdlg9OMgDiaxJRdQ365fpa+KGmhnYDSmI8VGzyGB+scCrsrocQj2+x2q
2Nk+/67TX6usUDZB1KVRutVrp/btJzbgT9qyCG6OMUse4hIPSAQ2BsMYcBo89tT2/x7HaN08iZlB
h1u5AlqlCp5yZZ/wRqcXzrdPrkyyezwA9+DOn1gwii+qCELuhbQOreCqZMV7utO2UXzA3k+LR5hh
bhQ/t93z+PKFxr/wFiROJYNhOCXxKCprgva6ALBaqI9XYe3OVa0SQfS7/ASHcWqhPMNJ+5IN/yFZ
kEZS1/vuw6mf+fkXrBI+7qLhc3Fj+CHfDSeN5sD4zAVe8cwBlE0G2Pl4oETXdBQt5CxyUEzZ+WQn
yKQggj9O58mxi3ZP9uou4UN6nBRS9xsHkrvbDSJ4e+Y8CuJ7/6a4I/l/EyuT/wxUfVBDKM5Dihm0
Ejw5c9nW4DZW/erpcV/VEB/eHsBQR78gGnq3u1PnxQrWNw9ZtjtdgPjRqnkUUtewi0Jpu4G9mTE1
0b/czGQVxG9AkjmRV/Vk1mutdKToLGhi4uAkjnIS8d6QXlZa+apWlUc8w4a5SFLsOB1qhrDVP0SF
EcK2RpqRQgvDLl2L1NLSCRMVF4VXQJ0LWu7c7qsKYU8VGDnNT9/fDLJyjliZxO+Dq9A58646qEvv
bqpYg0ArAxCsCYfFAz+9M76srGoCEmaUCnNkz48xJm+k2y6DqYc4V99iqa1saUFxYK7Qff1s0g7i
sNXLD8u5EJnzr9RS8ZsoVsc9vwufK32gmUmEoHJti+IW4gobWlSeItqZ6dTfX01KUTHzMIDQEbfy
nKOtzt3Ix2EcKmN/bAUHpD/QYTDaj0duOFdnq4mbUkHG/jaf1zBFMiUaEszbdXNKsoOmYR1jit3Z
aLh4+12YCXqNk5Sp9BPYxs8K+Iq/fZvWJdwRXNxxZMiQYaqYCoM0evm+oMjlmKKAQmBRuWXAqyho
+6Il9EgX3G9+8VKJHmwNcf1NkheUsgfDlVMBggxR7LeyW7TUrLLdCoEMXP7EwWYkvXpaEvHd71th
mgbP2QIbpw2z3//nWjPpEXH9lx92ixY0HUg2TcwKkdCAx5t0cOuP+1j6akmoEeEtHe2QXdDHeFxy
Yv1MSPbrlTH2coLDMfTUqC68ubtOly6CC9yNVTs6cTh2oDaTOs4iOCVrqpRV3KX8iOvtAd84HshH
s0Wf8+wfLVcQM9V7OMEt/DriHKGanHrOXHa32pzNetYi8zzWx+Sli/0GjvkxZanqdQ5OBPs4U09u
39+o51zekSg8MoaqeTbtC+1vdkNQcSYxTRHssG2xlLzZE1UAPqctuxvHo8LSGzBgISZgdbRHB4q3
SIQgvg/nJyAPwm1vMPnR6MWeL93hx1KOEu/bqVjGi84FCf8Fhx3gBaN/1suIkP/6rDiQ9oR5lId8
gPn1SscjPZoXTrXlujS9GHqGvNRUh+8PSnolDAPC6BtOZyPkTfFm80Mq22yMRRDUgy7Jwg55P+E9
DRF5zqRI395cvo6+sYX57a8ZXwHhCtpprwMd81JF+RBTfKq5TGYnFi/WU5WHUk4OcQXaPwt5WyXy
f6CwKXavbN25hWzv5o0ufSV5xK9IlutEhwHt5IXIO5VQg8za8UO2YpzZpmtP0ijfOzb9lHRB/7KP
6YEibCNZWMgORS6OE1FhCMR/rVR+M7h2RHYeK3vARFmoGvY/FUtjkg4H8kaC7VvlP5u6N1Sf+LZG
6BW1uw/WbZ7d8+o+9cWBXJcC7F22VW1DVbTFaRkfVvujIiuevjCEj8WTnY0rpltaO2AYaZc9qH2V
/EAK63Gd1siIhASXvP1jHpv2xwaUeRpcJpubA1w/LoxHkP3SIbHIyV93M2gGqAv3qU16ljQ9wWLk
bZG+QTT+F9u6ObgA5WgKWAUdY4OWfQ0Ut3gedEsRdKn22o/I/8S65+Mw6Xgpk+I2jV+8pzUa0UqF
rX4d/3Dtx7HNfzNweOvsaatQMHw2ueFIB308V6s0uAD4uzY0YsbWURKiMH1zRVQKaTiweOiZorDf
9vEVDvor9IUZoMBBkTcYrMBrWrgAJ5qz/h6DK2nH+mjP4uTJSTUSy+Hv6PMOtfn5l8JssygKdqiN
r5lqTBNMFTdoZugqSV3Wuu6/JXIPabDWiw==
`protect end_protected
